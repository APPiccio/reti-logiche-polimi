library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity project_tb is
end project_tb;
architecture projecttb of project_tb is
constant c_CLOCK_PERIOD		: time := 15 ns;
signal   tb_done		: std_logic;
signal   mem_address		: std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst		    : std_logic := '0';
signal   tb_start		: std_logic := '0';
signal   tb_clk		    : std_logic := '0';
signal   mem_o_data,mem_i_data		: std_logic_vector (7 downto 0);
signal   enable_wire  		: std_logic;
signal   mem_we		: std_logic;
type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
signal RAM: ram_type := (2 => "01010011", 3 => "00110011", 4 => "11000100",
 5 => "10011100",
 6 => "10001011",
 7 => "01000000",
 8 => "10010010",
 9 => "01010111",
 10 => "00110010",
 11 => "10010111",
 12 => "10101001",
 13 => "01000111",
 14 => "11110001",
 15 => "11101101",
 16 => "10111100",
 17 => "00001101",
 18 => "10001000",
 19 => "00110101",
 20 => "01110100",
 21 => "00011000",
 22 => "10000000",
 23 => "10011101",
 24 => "10100111",
 25 => "10101000",
 26 => "01010010",
 27 => "01110011",
 28 => "01000010",
 29 => "00101100",
 30 => "00000100",
 31 => "11001000",
 32 => "11110110",
 33 => "11000010",
 34 => "01000110",
 35 => "00000111",
 36 => "11110111",
 37 => "01010111",
 38 => "10000101",
 39 => "00011100",
 40 => "01100111",
 41 => "00011110",
 42 => "00101000",
 43 => "00110101",
 44 => "01000011",
 45 => "00011010",
 46 => "01001101",
 47 => "00111011",
 48 => "01011011",
 49 => "01111010",
 50 => "01010000",
 51 => "01101010",
 52 => "01000010",
 53 => "00110100",
 54 => "10011111",
 55 => "11111010",
 56 => "11011101",
 57 => "00100000",
 58 => "00101011",
 59 => "00111101",
 60 => "11001111",
 61 => "01010011",
 62 => "01010111",
 63 => "11001101",
 64 => "11000000",
 65 => "10100010",
 66 => "10000100",
 67 => "10011101",
 68 => "11100001",
 69 => "10101000",
 70 => "00101101",
 71 => "01000001",
 72 => "11110101",
 73 => "11001001",
 74 => "00001111",
 75 => "11001110",
 76 => "01001001",
 77 => "11001001",
 78 => "00101000",
 79 => "10110001",
 80 => "11011111",
 81 => "01000010",
 82 => "10000101",
 83 => "11110010",
 84 => "01100101",
 85 => "10011010",
 86 => "00110110",
 87 => "00011110",
 88 => "01010010",
 89 => "00000011",
 90 => "01010111",
 91 => "10010100",
 92 => "01100011",
 93 => "01001001",
 94 => "01110000",
 95 => "11110111",
 96 => "10111111",
 97 => "10101111",
 98 => "10001010",
 99 => "10011110",
 100 => "11101110",
 101 => "10101110",
 102 => "10111101",
 103 => "10111000",
 104 => "01001101",
 105 => "01001010",
 106 => "10000010",
 107 => "01000111",
 108 => "00000101",
 109 => "00000100",
 110 => "11010011",
 111 => "00010111",
 112 => "00010010",
 113 => "10001100",
 114 => "01100101",
 115 => "11111010",
 116 => "10101101",
 117 => "10110010",
 118 => "01011100",
 119 => "10100100",
 120 => "00010010",
 121 => "11100100",
 122 => "01101010",
 123 => "01100011",
 124 => "10000010",
 125 => "00011001",
 126 => "11110110",
 127 => "01111010",
 128 => "01010110",
 129 => "00001010",
 130 => "01100101",
 131 => "11011010",
 132 => "11110111",
 133 => "00101110",
 134 => "01110110",
 135 => "00101010",
 136 => "01011010",
 137 => "10001010",
 138 => "00110000",
 139 => "00010010",
 140 => "10111010",
 141 => "10111010",
 142 => "11110110",
 143 => "00010110",
 144 => "11011100",
 145 => "10010000",
 146 => "11111011",
 147 => "01101011",
 148 => "01001001",
 149 => "00110010",
 150 => "01011100",
 151 => "00000110",
 152 => "01111011",
 153 => "11011111",
 154 => "10010111",
 155 => "11001100",
 156 => "00010001",
 157 => "01011101",
 158 => "00000011",
 159 => "00000100",
 160 => "01110110",
 161 => "10000010",
 162 => "10001100",
 163 => "01101100",
 164 => "01101100",
 165 => "10000111",
 166 => "11000000",
 167 => "00101101",
 168 => "01111100",
 169 => "11001101",
 170 => "00001110",
 171 => "11000101",
 172 => "00000110",
 173 => "11110001",
 174 => "11110001",
 175 => "11101000",
 176 => "00010110",
 177 => "10100110",
 178 => "00101111",
 179 => "01110011",
 180 => "10100110",
 181 => "11111000",
 182 => "00101101",
 183 => "00010110",
 184 => "01000110",
 185 => "11000100",
 186 => "00101011",
 187 => "00010011",
 188 => "10010101",
 189 => "00001100",
 190 => "01111001",
 191 => "11000000",
 192 => "00110000",
 193 => "10111010",
 194 => "11100000",
 195 => "11100011",
 196 => "01001000",
 197 => "01101010",
 198 => "01111111",
 199 => "10110000",
 200 => "11111110",
 201 => "10011000",
 202 => "10111101",
 203 => "00110000",
 204 => "01101100",
 205 => "11011000",
 206 => "01100010",
 207 => "10001010",
 208 => "11110110",
 209 => "11010101",
 210 => "11010001",
 211 => "00110110",
 212 => "00000100",
 213 => "10000111",
 214 => "11111000",
 215 => "10011110",
 216 => "00000001",
 217 => "10010000",
 218 => "00101010",
 219 => "10111100",
 220 => "00001110",
 221 => "00011101",
 222 => "11100101",
 223 => "00111000",
 224 => "10111111",
 225 => "10000000",
 226 => "11101011",
 227 => "11010000",
 228 => "11001000",
 229 => "10000111",
 230 => "10001100",
 231 => "11001101",
 232 => "00011010",
 233 => "11100010",
 234 => "00101001",
 235 => "00001101",
 236 => "11101001",
 237 => "11100111",
 238 => "10101111",
 239 => "11000000",
 240 => "01111111",
 241 => "01110001",
 242 => "10100010",
 243 => "00011100",
 244 => "01000010",
 245 => "00100110",
 246 => "11010001",
 247 => "11000111",
 248 => "10110101",
 249 => "11111101",
 250 => "10101111",
 251 => "00111011",
 252 => "11011110",
 253 => "10100001",
 254 => "10010110",
 255 => "11001000",
 256 => "00011110",
 257 => "01100100",
 258 => "11111111",
 259 => "01101011",
 260 => "01101100",
 261 => "11111000",
 262 => "11010000",
 263 => "10010100",
 264 => "11101001",
 265 => "00010110",
 266 => "00000110",
 267 => "10100000",
 268 => "00010000",
 269 => "11001010",
 270 => "11001111",
 271 => "00101111",
 272 => "10011111",
 273 => "00101001",
 274 => "01000000",
 275 => "01101011",
 276 => "01011001",
 277 => "01001110",
 278 => "01100010",
 279 => "00101001",
 280 => "00001011",
 281 => "11001111",
 282 => "01111000",
 283 => "01000101",
 284 => "01111100",
 285 => "10010110",
 286 => "10101111",
 287 => "10011100",
 288 => "10110111",
 289 => "01101010",
 290 => "00010110",
 291 => "01111011",
 292 => "10000011",
 293 => "01001111",
 294 => "11011011",
 295 => "10101010",
 296 => "10000100",
 297 => "00011001",
 298 => "01000011",
 299 => "11010101",
 300 => "11000111",
 301 => "01101011",
 302 => "11001011",
 303 => "11011101",
 304 => "10011011",
 305 => "10101010",
 306 => "10000010",
 307 => "10100101",
 308 => "00111110",
 309 => "01000101",
 310 => "00001110",
 311 => "11001110",
 312 => "11000000",
 313 => "10001111",
 314 => "11010000",
 315 => "01110010",
 316 => "11010111",
 317 => "10001011",
 318 => "00001101",
 319 => "00010000",
 320 => "01011001",
 321 => "11011001",
 322 => "01000101",
 323 => "10111100",
 324 => "11001111",
 325 => "00100111",
 326 => "11100100",
 327 => "10111110",
 328 => "10011001",
 329 => "10000010",
 330 => "11010111",
 331 => "11001111",
 332 => "10110100",
 333 => "00101110",
 334 => "01100000",
 335 => "10101000",
 336 => "00110101",
 337 => "01101101",
 338 => "01100011",
 339 => "00001110",
 340 => "10001000",
 341 => "10111001",
 342 => "01100100",
 343 => "00001011",
 344 => "11010010",
 345 => "11100101",
 346 => "00000100",
 347 => "11100010",
 348 => "11010001",
 349 => "00100101",
 350 => "10001100",
 351 => "10110000",
 352 => "11100011",
 353 => "10011010",
 354 => "00010101",
 355 => "11001111",
 356 => "11100010",
 357 => "10000111",
 358 => "01010101",
 359 => "00010110",
 360 => "10100000",
 361 => "11001111",
 362 => "00001101",
 363 => "00011001",
 364 => "01110100",
 365 => "01010011",
 366 => "11110000",
 367 => "11000010",
 368 => "11101001",
 369 => "11110111",
 370 => "00011010",
 371 => "11000000",
 372 => "00011010",
 373 => "01100000",
 374 => "11010101",
 375 => "00001110",
 376 => "00111010",
 377 => "11110101",
 378 => "11110001",
 379 => "00000001",
 380 => "00001100",
 381 => "10101101",
 382 => "00000111",
 383 => "00000001",
 384 => "10011110",
 385 => "11010110",
 386 => "10001010",
 387 => "01110000",
 388 => "01100010",
 389 => "01110001",
 390 => "11000100",
 391 => "10110110",
 392 => "00000000",
 393 => "00101011",
 394 => "00111101",
 395 => "11111000",
 396 => "01111110",
 397 => "11100001",
 398 => "01001010",
 399 => "10111111",
 400 => "01001111",
 401 => "10101110",
 402 => "01100000",
 403 => "11110110",
 404 => "10001000",
 405 => "00010110",
 406 => "10100000",
 407 => "11111001",
 408 => "10010100",
 409 => "00101011",
 410 => "11010010",
 411 => "00010100",
 412 => "10011000",
 413 => "01110001",
 414 => "00001100",
 415 => "01100010",
 416 => "00111110",
 417 => "01101100",
 418 => "10011110",
 419 => "11011111",
 420 => "11001100",
 421 => "00111000",
 422 => "00110111",
 423 => "01001000",
 424 => "10010011",
 425 => "11001010",
 426 => "10011110",
 427 => "00000000",
 428 => "10110110",
 429 => "10010101",
 430 => "11011100",
 431 => "00110100",
 432 => "01011100",
 433 => "11110010",
 434 => "01010100",
 435 => "10101011",
 436 => "01000011",
 437 => "01010100",
 438 => "00000011",
 439 => "10101100",
 440 => "10100010",
 441 => "01010011",
 442 => "01101100",
 443 => "01101000",
 444 => "01111000",
 445 => "01010111",
 446 => "11101001",
 447 => "01110001",
 448 => "00100101",
 449 => "00011101",
 450 => "00110111",
 451 => "11100100",
 452 => "10110100",
 453 => "00010101",
 454 => "01100000",
 455 => "11000100",
 456 => "01000101",
 457 => "00000001",
 458 => "01000010",
 459 => "11011110",
 460 => "11001101",
 461 => "11111110",
 462 => "10101110",
 463 => "10001100",
 464 => "01101111",
 465 => "00110101",
 466 => "01110100",
 467 => "00001010",
 468 => "11011100",
 469 => "00011000",
 470 => "11010001",
 471 => "01110100",
 472 => "10111110",
 473 => "00110010",
 474 => "01010110",
 475 => "01000111",
 476 => "00111010",
 477 => "10001111",
 478 => "00100111",
 479 => "11110000",
 480 => "01000000",
 481 => "00111110",
 482 => "00000011",
 483 => "10101101",
 484 => "00100000",
 485 => "11100111",
 486 => "00001101",
 487 => "01001101",
 488 => "10001011",
 489 => "10111100",
 490 => "10100000",
 491 => "01101010",
 492 => "10010010",
 493 => "10100010",
 494 => "10001010",
 495 => "01011001",
 496 => "10110110",
 497 => "00101101",
 498 => "00010100",
 499 => "10000101",
 500 => "10000000",
 501 => "01111000",
 502 => "11010110",
 503 => "11011010",
 504 => "01011011",
 505 => "11111010",
 506 => "10100011",
 507 => "00110000",
 508 => "10001000",
 509 => "00000100",
 510 => "01110001",
 511 => "01000100",
 512 => "00101001",
 513 => "00100111",
 514 => "10101111",
 515 => "10010100",
 516 => "00000001",
 517 => "11000010",
 518 => "00000001",
 519 => "10110100",
 520 => "00010101",
 521 => "11010010",
 522 => "11000000",
 523 => "00011110",
 524 => "00011000",
 525 => "10001000",
 526 => "10111010",
 527 => "11101101",
 528 => "10000100",
 529 => "10001000",
 530 => "01101101",
 531 => "01001011",
 532 => "10000010",
 533 => "10011100",
 534 => "11010011",
 535 => "10010101",
 536 => "10011110",
 537 => "00111010",
 538 => "11001101",
 539 => "01100100",
 540 => "10111000",
 541 => "10101001",
 542 => "00100101",
 543 => "10010000",
 544 => "00000011",
 545 => "00110000",
 546 => "11010111",
 547 => "11110111",
 548 => "00101011",
 549 => "01001000",
 550 => "11000111",
 551 => "11101001",
 552 => "11110111",
 553 => "10100100",
 554 => "10000111",
 555 => "11100011",
 556 => "00100101",
 557 => "00110110",
 558 => "00011000",
 559 => "01101001",
 560 => "10101100",
 561 => "11100111",
 562 => "11110011",
 563 => "10100100",
 564 => "10010101",
 565 => "11000010",
 566 => "00000110",
 567 => "00100000",
 568 => "00110111",
 569 => "11110010",
 570 => "10101000",
 571 => "11001100",
 572 => "10110101",
 573 => "11100100",
 574 => "11001010",
 575 => "10101001",
 576 => "11101010",
 577 => "10110111",
 578 => "01000100",
 579 => "10001010",
 580 => "11000010",
 581 => "10010010",
 582 => "01110111",
 583 => "01111000",
 584 => "11000100",
 585 => "01110101",
 586 => "00010001",
 587 => "10001011",
 588 => "01100010",
 589 => "00110001",
 590 => "01011000",
 591 => "10101100",
 592 => "11111100",
 593 => "00110100",
 594 => "10010000",
 595 => "00001100",
 596 => "00101111",
 597 => "10110110",
 598 => "00001000",
 599 => "11000001",
 600 => "11011100",
 601 => "11111101",
 602 => "10100001",
 603 => "01111001",
 604 => "00001010",
 605 => "11000101",
 606 => "10001000",
 607 => "11101011",
 608 => "11010111",
 609 => "10100010",
 610 => "00001011",
 611 => "00010000",
 612 => "00010000",
 613 => "00010110",
 614 => "11000000",
 615 => "00011011",
 616 => "11100010",
 617 => "11011110",
 618 => "10110001",
 619 => "01101111",
 620 => "00001111",
 621 => "10100111",
 622 => "10001010",
 623 => "10100001",
 624 => "01101101",
 625 => "11010100",
 626 => "00010010",
 627 => "01011100",
 628 => "01100110",
 629 => "10100101",
 630 => "01101001",
 631 => "10011001",
 632 => "00111110",
 633 => "01011110",
 634 => "01010010",
 635 => "11101110",
 636 => "01011010",
 637 => "00100111",
 638 => "11001101",
 639 => "00001011",
 640 => "10010101",
 641 => "00010101",
 642 => "10001000",
 643 => "10111010",
 644 => "10111110",
 645 => "11101011",
 646 => "01110000",
 647 => "10110100",
 648 => "01110010",
 649 => "11111011",
 650 => "00111101",
 651 => "00111010",
 652 => "10111010",
 653 => "11000110",
 654 => "00101000",
 655 => "11101110",
 656 => "01100111",
 657 => "00111100",
 658 => "11101001",
 659 => "11100111",
 660 => "00110101",
 661 => "11000111",
 662 => "00011000",
 663 => "10101010",
 664 => "01111000",
 665 => "01000111",
 666 => "00101110",
 667 => "10101100",
 668 => "11000000",
 669 => "01110010",
 670 => "10111001",
 671 => "11011001",
 672 => "11000001",
 673 => "10101101",
 674 => "11010110",
 675 => "10000000",
 676 => "00000101",
 677 => "00111110",
 678 => "10011101",
 679 => "00110100",
 680 => "10010010",
 681 => "00011011",
 682 => "01100001",
 683 => "10111110",
 684 => "11111010",
 685 => "01111110",
 686 => "00111101",
 687 => "00110001",
 688 => "01000101",
 689 => "00001000",
 690 => "01011000",
 691 => "00110001",
 692 => "00000111",
 693 => "00010000",
 694 => "11100100",
 695 => "11110100",
 696 => "10000000",
 697 => "01111111",
 698 => "10010101",
 699 => "11100010",
 700 => "10010010",
 701 => "01001101",
 702 => "11011101",
 703 => "01001110",
 704 => "00100000",
 705 => "01101110",
 706 => "10101010",
 707 => "01101100",
 708 => "01101001",
 709 => "01011110",
 710 => "00010110",
 711 => "00001011",
 712 => "11100001",
 713 => "11110111",
 714 => "01000100",
 715 => "11001100",
 716 => "10111101",
 717 => "11110010",
 718 => "01100111",
 719 => "11100110",
 720 => "11010011",
 721 => "00011010",
 722 => "01100110",
 723 => "11110110",
 724 => "10111011",
 725 => "00000100",
 726 => "11011011",
 727 => "00000001",
 728 => "10110010",
 729 => "00011000",
 730 => "10000100",
 731 => "10011010",
 732 => "11000100",
 733 => "11010101",
 734 => "01100100",
 735 => "00110101",
 736 => "10100101",
 737 => "01100000",
 738 => "11110101",
 739 => "00101101",
 740 => "00110011",
 741 => "11010001",
 742 => "01000111",
 743 => "10000111",
 744 => "11100101",
 745 => "11100011",
 746 => "10110001",
 747 => "01011000",
 748 => "11001111",
 749 => "01000010",
 750 => "00101001",
 751 => "01000011",
 752 => "00000111",
 753 => "11000100",
 754 => "10101000",
 755 => "01101000",
 756 => "10001011",
 757 => "11010100",
 758 => "00000110",
 759 => "10011001",
 760 => "11001100",
 761 => "11110010",
 762 => "00001111",
 763 => "00101010",
 764 => "11101100",
 765 => "11011111",
 766 => "11110010",
 767 => "10010010",
 768 => "01010100",
 769 => "11100110",
 770 => "10000101",
 771 => "01001011",
 772 => "11001011",
 773 => "11001000",
 774 => "10010000",
 775 => "10011001",
 776 => "00110001",
 777 => "10101011",
 778 => "00110010",
 779 => "11010010",
 780 => "00101010",
 781 => "00111100",
 782 => "10000110",
 783 => "10001111",
 784 => "10111111",
 785 => "01010101",
 786 => "00110110",
 787 => "11111100",
 788 => "01001000",
 789 => "10101101",
 790 => "11100011",
 791 => "10101101",
 792 => "10011001",
 793 => "11011010",
 794 => "11111000",
 795 => "01101010",
 796 => "01000000",
 797 => "01100110",
 798 => "10010111",
 799 => "00010100",
 800 => "00000001",
 801 => "01101011",
 802 => "01100001",
 803 => "01101110",
 804 => "00100000",
 805 => "00100001",
 806 => "00101001",
 807 => "01100000",
 808 => "01001001",
 809 => "10001001",
 810 => "11100000",
 811 => "01010010",
 812 => "10110000",
 813 => "10101111",
 814 => "00010011",
 815 => "00100001",
 816 => "11000001",
 817 => "11110110",
 818 => "10000110",
 819 => "11001011",
 820 => "10101110",
 821 => "01010001",
 822 => "11100101",
 823 => "01110011",
 824 => "10001011",
 825 => "10101001",
 826 => "00000001",
 827 => "11101000",
 828 => "10101100",
 829 => "10100000",
 830 => "10100100",
 831 => "11000011",
 832 => "00010101",
 833 => "11111010",
 834 => "01111110",
 835 => "11000011",
 836 => "00001001",
 837 => "11001111",
 838 => "00111100",
 839 => "00101110",
 840 => "00111011",
 841 => "01001110",
 842 => "00010010",
 843 => "01100111",
 844 => "00011111",
 845 => "10010101",
 846 => "01000000",
 847 => "01000010",
 848 => "11110001",
 849 => "11111110",
 850 => "00100010",
 851 => "00110011",
 852 => "00011011",
 853 => "00101110",
 854 => "10111111",
 855 => "00111110",
 856 => "11101010",
 857 => "01001100",
 858 => "11000001",
 859 => "00101101",
 860 => "00110001",
 861 => "00011000",
 862 => "00001011",
 863 => "10000110",
 864 => "00001101",
 865 => "10010111",
 866 => "10100011",
 867 => "00001110",
 868 => "11010001",
 869 => "01100001",
 870 => "00010111",
 871 => "00001011",
 872 => "11111000",
 873 => "11000101",
 874 => "11000000",
 875 => "10011011",
 876 => "00000001",
 877 => "11011001",
 878 => "01111100",
 879 => "00101001",
 880 => "10001001",
 881 => "00100100",
 882 => "00101111",
 883 => "10001010",
 884 => "10111100",
 885 => "00000011",
 886 => "01100111",
 887 => "00100010",
 888 => "11100110",
 889 => "01101010",
 890 => "11001101",
 891 => "11011110",
 892 => "11001001",
 893 => "10001001",
 894 => "11110010",
 895 => "10011110",
 896 => "00111010",
 897 => "10000010",
 898 => "01111001",
 899 => "00001000",
 900 => "10011011",
 901 => "00100011",
 902 => "00100100",
 903 => "11101100",
 904 => "11001110",
 905 => "10011110",
 906 => "00010011",
 907 => "11001101",
 908 => "10111111",
 909 => "10101000",
 910 => "10001000",
 911 => "10000110",
 912 => "01000010",
 913 => "01001010",
 914 => "10010000",
 915 => "00111011",
 916 => "01100111",
 917 => "10011011",
 918 => "00011010",
 919 => "01101010",
 920 => "01100011",
 921 => "00010111",
 922 => "01100000",
 923 => "01111110",
 924 => "10010101",
 925 => "11110111",
 926 => "00010110",
 927 => "11100101",
 928 => "10101011",
 929 => "00011101",
 930 => "11010000",
 931 => "01001110",
 932 => "00001101",
 933 => "10011001",
 934 => "00001010",
 935 => "11111110",
 936 => "11010101",
 937 => "10000111",
 938 => "00110101",
 939 => "10000000",
 940 => "00011000",
 941 => "11000010",
 942 => "01101001",
 943 => "00100000",
 944 => "01011010",
 945 => "11111100",
 946 => "00010111",
 947 => "11101100",
 948 => "10100001",
 949 => "10101110",
 950 => "00010110",
 951 => "11101010",
 952 => "10010010",
 953 => "10100001",
 954 => "01111111",
 955 => "11100111",
 956 => "11101011",
 957 => "11001111",
 958 => "00111001",
 959 => "10110010",
 960 => "01010101",
 961 => "00011111",
 962 => "00101100",
 963 => "01101010",
 964 => "00011101",
 965 => "00110111",
 966 => "01010001",
 967 => "00010101",
 968 => "11100000",
 969 => "11011111",
 970 => "11011011",
 971 => "10101010",
 972 => "11111010",
 973 => "00101010",
 974 => "11011111",
 975 => "00110011",
 976 => "00111110",
 977 => "11001111",
 978 => "01010100",
 979 => "10000001",
 980 => "10100110",
 981 => "11001100",
 982 => "10001100",
 983 => "00010110",
 984 => "11010101",
 985 => "11010000",
 986 => "10100001",
 987 => "11011011",
 988 => "11001000",
 989 => "11000101",
 990 => "11100011",
 991 => "01000101",
 992 => "10000001",
 993 => "10111000",
 994 => "10011111",
 995 => "00100000",
 996 => "10000101",
 997 => "01001101",
 998 => "00000111",
 999 => "11000110",
 1000 => "01100000",
 1001 => "10100010",
 1002 => "10001101",
 1003 => "10111010",
 1004 => "10101110",
 1005 => "01010100",
 1006 => "11101100",
 1007 => "10101111",
 1008 => "01000110",
 1009 => "10101110",
 1010 => "01011011",
 1011 => "00100011",
 1012 => "10111001",
 1013 => "00110010",
 1014 => "10010001",
 1015 => "01100110",
 1016 => "00110000",
 1017 => "11010101",
 1018 => "00011100",
 1019 => "11101100",
 1020 => "11011101",
 1021 => "11110011",
 1022 => "00000011",
 1023 => "11000101",
 1024 => "11010101",
 1025 => "10101111",
 1026 => "10111001",
 1027 => "01000001",
 1028 => "00011001",
 1029 => "11010000",
 1030 => "01101011",
 1031 => "00110000",
 1032 => "11110101",
 1033 => "10001101",
 1034 => "11010111",
 1035 => "01011011",
 1036 => "11001101",
 1037 => "11010001",
 1038 => "10001110",
 1039 => "00000110",
 1040 => "00001111",
 1041 => "00000110",
 1042 => "10001000",
 1043 => "11001011",
 1044 => "11100010",
 1045 => "10000001",
 1046 => "10011001",
 1047 => "10111000",
 1048 => "11111001",
 1049 => "00111011",
 1050 => "10110010",
 1051 => "01000001",
 1052 => "01101111",
 1053 => "11100011",
 1054 => "11111101",
 1055 => "11010110",
 1056 => "11001011",
 1057 => "10001011",
 1058 => "10110100",
 1059 => "10110111",
 1060 => "10010010",
 1061 => "11110010",
 1062 => "10100111",
 1063 => "00000100",
 1064 => "01000001",
 1065 => "00111011",
 1066 => "11000010",
 1067 => "10011000",
 1068 => "10100110",
 1069 => "11011111",
 1070 => "01011101",
 1071 => "01010110",
 1072 => "10011110",
 1073 => "11000101",
 1074 => "00001001",
 1075 => "00100110",
 1076 => "11011001",
 1077 => "00111100",
 1078 => "01001111",
 1079 => "00010100",
 1080 => "01001011",
 1081 => "01111001",
 1082 => "00110000",
 1083 => "11001001",
 1084 => "00100110",
 1085 => "01111111",
 1086 => "10001010",
 1087 => "01001001",
 1088 => "01010110",
 1089 => "01011101",
 1090 => "11110011",
 1091 => "00011001",
 1092 => "10010001",
 1093 => "01001011",
 1094 => "01101011",
 1095 => "11111110",
 1096 => "10100000",
 1097 => "10110111",
 1098 => "11001000",
 1099 => "00000011",
 1100 => "01011001",
 1101 => "10011010",
 1102 => "11111010",
 1103 => "00110000",
 1104 => "11000100",
 1105 => "01010101",
 1106 => "00011010",
 1107 => "01011101",
 1108 => "11100001",
 1109 => "10010110",
 1110 => "01000100",
 1111 => "10011011",
 1112 => "10100001",
 1113 => "00111101",
 1114 => "11011001",
 1115 => "01001101",
 1116 => "01000110",
 1117 => "11110101",
 1118 => "01111011",
 1119 => "00110111",
 1120 => "01000000",
 1121 => "01110110",
 1122 => "00010010",
 1123 => "10110001",
 1124 => "10000001",
 1125 => "10011001",
 1126 => "00110001",
 1127 => "11110010",
 1128 => "11000111",
 1129 => "11010100",
 1130 => "11100001",
 1131 => "11101100",
 1132 => "11011101",
 1133 => "01011110",
 1134 => "01100000",
 1135 => "01100001",
 1136 => "11001001",
 1137 => "00010001",
 1138 => "10101110",
 1139 => "00101011",
 1140 => "00110011",
 1141 => "00111001",
 1142 => "10011010",
 1143 => "11000001",
 1144 => "10100110",
 1145 => "11001111",
 1146 => "00010100",
 1147 => "10101011",
 1148 => "01010101",
 1149 => "10110101",
 1150 => "01111111",
 1151 => "10110110",
 1152 => "01101111",
 1153 => "10001000",
 1154 => "01100101",
 1155 => "01110010",
 1156 => "00010010",
 1157 => "01001111",
 1158 => "01101011",
 1159 => "11010011",
 1160 => "01000001",
 1161 => "00100011",
 1162 => "00110010",
 1163 => "10000001",
 1164 => "10010011",
 1165 => "01000101",
 1166 => "00110111",
 1167 => "11110111",
 1168 => "11111100",
 1169 => "01101111",
 1170 => "01110111",
 1171 => "11011100",
 1172 => "11111000",
 1173 => "11010111",
 1174 => "11000111",
 1175 => "00001000",
 1176 => "10100000",
 1177 => "11011100",
 1178 => "01000101",
 1179 => "11100011",
 1180 => "11001011",
 1181 => "01001010",
 1182 => "00000001",
 1183 => "11011110",
 1184 => "11000011",
 1185 => "11011010",
 1186 => "01011001",
 1187 => "00111001",
 1188 => "11101000",
 1189 => "01001100",
 1190 => "10101001",
 1191 => "01001011",
 1192 => "00111101",
 1193 => "01010001",
 1194 => "10000011",
 1195 => "01111101",
 1196 => "01001100",
 1197 => "00011001",
 1198 => "01101000",
 1199 => "11101111",
 1200 => "10111010",
 1201 => "01110101",
 1202 => "01111111",
 1203 => "01011010",
 1204 => "10101001",
 1205 => "00000011",
 1206 => "10111011",
 1207 => "00111011",
 1208 => "01010010",
 1209 => "10111010",
 1210 => "10101000",
 1211 => "01111100",
 1212 => "01011000",
 1213 => "10101011",
 1214 => "10100001",
 1215 => "00010100",
 1216 => "01011011",
 1217 => "10100111",
 1218 => "01100110",
 1219 => "10111011",
 1220 => "01000011",
 1221 => "00100110",
 1222 => "01011010",
 1223 => "01001011",
 1224 => "00100001",
 1225 => "01101100",
 1226 => "10001001",
 1227 => "01001110",
 1228 => "01110111",
 1229 => "11010101",
 1230 => "10011100",
 1231 => "10110110",
 1232 => "01111000",
 1233 => "11011010",
 1234 => "01101101",
 1235 => "11100000",
 1236 => "11110001",
 1237 => "00111100",
 1238 => "01010000",
 1239 => "10001001",
 1240 => "11010011",
 1241 => "01000001",
 1242 => "01000100",
 1243 => "10011011",
 1244 => "01000110",
 1245 => "11011001",
 1246 => "10010110",
 1247 => "00001110",
 1248 => "00110000",
 1249 => "01001110",
 1250 => "01111000",
 1251 => "01010000",
 1252 => "11111011",
 1253 => "00110001",
 1254 => "10001000",
 1255 => "11111000",
 1256 => "01110100",
 1257 => "11111110",
 1258 => "01000100",
 1259 => "01111101",
 1260 => "11001001",
 1261 => "10011111",
 1262 => "00011111",
 1263 => "00111111",
 1264 => "10100010",
 1265 => "00110011",
 1266 => "01000101",
 1267 => "10100001",
 1268 => "00000101",
 1269 => "00001110",
 1270 => "11101000",
 1271 => "01010000",
 1272 => "01001101",
 1273 => "00111100",
 1274 => "00101010",
 1275 => "10001110",
 1276 => "11101011",
 1277 => "11100100",
 1278 => "10001010",
 1279 => "11010111",
 1280 => "10001110",
 1281 => "10100010",
 1282 => "01111100",
 1283 => "01100101",
 1284 => "11010011",
 1285 => "11101011",
 1286 => "01110111",
 1287 => "01110010",
 1288 => "10101110",
 1289 => "10001011",
 1290 => "01010100",
 1291 => "11100000",
 1292 => "11010101",
 1293 => "11001011",
 1294 => "11101010",
 1295 => "11100001",
 1296 => "01111110",
 1297 => "00110001",
 1298 => "01101100",
 1299 => "10110101",
 1300 => "00110010",
 1301 => "10000000",
 1302 => "10000100",
 1303 => "11111101",
 1304 => "01111001",
 1305 => "01110111",
 1306 => "10110011",
 1307 => "11001011",
 1308 => "11010000",
 1309 => "10101100",
 1310 => "00101111",
 1311 => "10110011",
 1312 => "01111111",
 1313 => "11000000",
 1314 => "10011110",
 1315 => "00001000",
 1316 => "10110111",
 1317 => "00000100",
 1318 => "00100010",
 1319 => "10101100",
 1320 => "00011110",
 1321 => "01100110",
 1322 => "01010110",
 1323 => "01001111",
 1324 => "01100100",
 1325 => "00001001",
 1326 => "00111010",
 1327 => "11001001",
 1328 => "00111010",
 1329 => "10100000",
 1330 => "00011010",
 1331 => "10101000",
 1332 => "10111011",
 1333 => "01110010",
 1334 => "01001100",
 1335 => "10010100",
 1336 => "11011100",
 1337 => "11100001",
 1338 => "10001011",
 1339 => "00011111",
 1340 => "00101110",
 1341 => "10100111",
 1342 => "01010000",
 1343 => "11101111",
 1344 => "00011000",
 1345 => "11110100",
 1346 => "01010111",
 1347 => "10110100",
 1348 => "01101010",
 1349 => "11101101",
 1350 => "01001111",
 1351 => "01101011",
 1352 => "00111111",
 1353 => "10110100",
 1354 => "10101001",
 1355 => "11110000",
 1356 => "10111101",
 1357 => "00110110",
 1358 => "01000011",
 1359 => "11100101",
 1360 => "00111101",
 1361 => "10111010",
 1362 => "01110100",
 1363 => "10100001",
 1364 => "01110011",
 1365 => "00010011",
 1366 => "00110001",
 1367 => "11100000",
 1368 => "10100110",
 1369 => "10100100",
 1370 => "10010100",
 1371 => "00010101",
 1372 => "10001000",
 1373 => "01100100",
 1374 => "01110100",
 1375 => "11111100",
 1376 => "00001000",
 1377 => "11111101",
 1378 => "10000001",
 1379 => "10100000",
 1380 => "11011110",
 1381 => "10111100",
 1382 => "10011110",
 1383 => "00011100",
 1384 => "10100110",
 1385 => "11101010",
 1386 => "01100100",
 1387 => "01100001",
 1388 => "10011001",
 1389 => "11010100",
 1390 => "11101010",
 1391 => "00001001",
 1392 => "10001011",
 1393 => "01111110",
 1394 => "11101101",
 1395 => "00101111",
 1396 => "01111100",
 1397 => "00011100",
 1398 => "00111011",
 1399 => "00000111",
 1400 => "11110000",
 1401 => "01011101",
 1402 => "11001111",
 1403 => "10010000",
 1404 => "00111101",
 1405 => "01101000",
 1406 => "01110111",
 1407 => "00111001",
 1408 => "11011111",
 1409 => "00011101",
 1410 => "11100001",
 1411 => "11100000",
 1412 => "00000111",
 1413 => "10101000",
 1414 => "01010011",
 1415 => "11100111",
 1416 => "01101101",
 1417 => "01010011",
 1418 => "00001111",
 1419 => "11100101",
 1420 => "01110010",
 1421 => "00100000",
 1422 => "11111101",
 1423 => "00010001",
 1424 => "00101011",
 1425 => "00110100",
 1426 => "11010101",
 1427 => "01001100",
 1428 => "00011000",
 1429 => "10111101",
 1430 => "00111011",
 1431 => "01111110",
 1432 => "11011011",
 1433 => "00011010",
 1434 => "01001111",
 1435 => "01000111",
 1436 => "10100000",
 1437 => "10001011",
 1438 => "00110001",
 1439 => "01011011",
 1440 => "11001000",
 1441 => "01010110",
 1442 => "00101001",
 1443 => "10100000",
 1444 => "11100110",
 1445 => "10000100",
 1446 => "00001001",
 1447 => "11110101",
 1448 => "11111101",
 1449 => "00111101",
 1450 => "10101101",
 1451 => "10001011",
 1452 => "00001111",
 1453 => "00000000",
 1454 => "10000100",
 1455 => "10001111",
 1456 => "11011000",
 1457 => "11001010",
 1458 => "10001011",
 1459 => "01001011",
 1460 => "01001011",
 1461 => "10000011",
 1462 => "01010100",
 1463 => "10110001",
 1464 => "11010010",
 1465 => "00010011",
 1466 => "00101110",
 1467 => "11100111",
 1468 => "01110011",
 1469 => "01010011",
 1470 => "10111010",
 1471 => "01010110",
 1472 => "10111100",
 1473 => "00000011",
 1474 => "11010100",
 1475 => "11001101",
 1476 => "11100001",
 1477 => "10101100",
 1478 => "00110101",
 1479 => "01101010",
 1480 => "01101111",
 1481 => "10001011",
 1482 => "10110101",
 1483 => "11110110",
 1484 => "10001110",
 1485 => "10010000",
 1486 => "00111010",
 1487 => "00111000",
 1488 => "10011000",
 1489 => "10100011",
 1490 => "11001111",
 1491 => "00100101",
 1492 => "00001110",
 1493 => "11011001",
 1494 => "01101001",
 1495 => "10010000",
 1496 => "11000101",
 1497 => "10100111",
 1498 => "00011101",
 1499 => "01110100",
 1500 => "01100000",
 1501 => "00010010",
 1502 => "00001000",
 1503 => "00000111",
 1504 => "01010011",
 1505 => "10011011",
 1506 => "01100101",
 1507 => "10110101",
 1508 => "10101001",
 1509 => "10011011",
 1510 => "10101110",
 1511 => "01100110",
 1512 => "10111011",
 1513 => "11100111",
 1514 => "11110001",
 1515 => "01011000",
 1516 => "00111000",
 1517 => "10100000",
 1518 => "10110000",
 1519 => "11001111",
 1520 => "01111110",
 1521 => "10011010",
 1522 => "11111111",
 1523 => "01000000",
 1524 => "10011000",
 1525 => "11101011",
 1526 => "01101101",
 1527 => "00110100",
 1528 => "10000011",
 1529 => "11000110",
 1530 => "11010110",
 1531 => "01000111",
 1532 => "10000110",
 1533 => "00100111",
 1534 => "10101110",
 1535 => "10010100",
 1536 => "00111110",
 1537 => "11011101",
 1538 => "10100010",
 1539 => "10010110",
 1540 => "00101111",
 1541 => "01111011",
 1542 => "00110111",
 1543 => "10000110",
 1544 => "10100100",
 1545 => "11110010",
 1546 => "01110010",
 1547 => "11010001",
 1548 => "10110100",
 1549 => "10110001",
 1550 => "00010101",
 1551 => "10111110",
 1552 => "00100100",
 1553 => "11111010",
 1554 => "11001110",
 1555 => "10011101",
 1556 => "00011111",
 1557 => "00000110",
 1558 => "11101100",
 1559 => "00101011",
 1560 => "01000001",
 1561 => "10001110",
 1562 => "11001000",
 1563 => "10111001",
 1564 => "00011101",
 1565 => "11001101",
 1566 => "01001100",
 1567 => "11011111",
 1568 => "01010101",
 1569 => "01111111",
 1570 => "01000000",
 1571 => "10100110",
 1572 => "10010101",
 1573 => "00001010",
 1574 => "01101101",
 1575 => "11000001",
 1576 => "11111001",
 1577 => "10011000",
 1578 => "11001011",
 1579 => "10111100",
 1580 => "01101011",
 1581 => "00111111",
 1582 => "11110110",
 1583 => "11111100",
 1584 => "10111111",
 1585 => "11111100",
 1586 => "11110011",
 1587 => "11100111",
 1588 => "00111010",
 1589 => "10100001",
 1590 => "00000100",
 1591 => "01011010",
 1592 => "11111000",
 1593 => "00100100",
 1594 => "00111000",
 1595 => "11001101",
 1596 => "10010011",
 1597 => "10001110",
 1598 => "01011011",
 1599 => "10011001",
 1600 => "11111001",
 1601 => "10001111",
 1602 => "00110011",
 1603 => "00110100",
 1604 => "00100100",
 1605 => "11100010",
 1606 => "00010101",
 1607 => "00100110",
 1608 => "11010100",
 1609 => "00010110",
 1610 => "00100100",
 1611 => "00011111",
 1612 => "01111110",
 1613 => "01111111",
 1614 => "01100100",
 1615 => "00000111",
 1616 => "01000001",
 1617 => "10110010",
 1618 => "10101101",
 1619 => "11101010",
 1620 => "00010001",
 1621 => "01010010",
 1622 => "10101000",
 1623 => "00010010",
 1624 => "10100110",
 1625 => "00111000",
 1626 => "10100000",
 1627 => "01010001",
 1628 => "00001110",
 1629 => "10010110",
 1630 => "11101001",
 1631 => "01010000",
 1632 => "01000010",
 1633 => "01011110",
 1634 => "10101001",
 1635 => "10110111",
 1636 => "01101001",
 1637 => "10010011",
 1638 => "01111011",
 1639 => "11001111",
 1640 => "11100000",
 1641 => "00101001",
 1642 => "11100100",
 1643 => "01101111",
 1644 => "00101000",
 1645 => "01101000",
 1646 => "11101000",
 1647 => "11111011",
 1648 => "00110110",
 1649 => "00111011",
 1650 => "01100100",
 1651 => "11111100",
 1652 => "00111001",
 1653 => "00110000",
 1654 => "00101010",
 1655 => "00001110",
 1656 => "00001001",
 1657 => "01110110",
 1658 => "01100011",
 1659 => "10011000",
 1660 => "10011110",
 1661 => "10001100",
 1662 => "10010001",
 1663 => "01010010",
 1664 => "10100101",
 1665 => "01101010",
 1666 => "10111100",
 1667 => "00000001",
 1668 => "00011100",
 1669 => "01111011",
 1670 => "10011100",
 1671 => "00001101",
 1672 => "01101111",
 1673 => "10101110",
 1674 => "11110010",
 1675 => "10000010",
 1676 => "10111010",
 1677 => "00100001",
 1678 => "01000110",
 1679 => "00111011",
 1680 => "11001011",
 1681 => "01001101",
 1682 => "11111010",
 1683 => "01011111",
 1684 => "01001101",
 1685 => "00101100",
 1686 => "10001000",
 1687 => "11011011",
 1688 => "00100111",
 1689 => "10011110",
 1690 => "11101110",
 1691 => "11101011",
 1692 => "11100101",
 1693 => "10010101",
 1694 => "01010100",
 1695 => "01101000",
 1696 => "00001011",
 1697 => "10100100",
 1698 => "11011111",
 1699 => "00011111",
 1700 => "10110111",
 1701 => "00001111",
 1702 => "00011000",
 1703 => "11101001",
 1704 => "10000000",
 1705 => "10010110",
 1706 => "11001100",
 1707 => "11111000",
 1708 => "11100001",
 1709 => "10100100",
 1710 => "01100110",
 1711 => "11001010",
 1712 => "01101111",
 1713 => "10110001",
 1714 => "01100101",
 1715 => "11001110",
 1716 => "11001010",
 1717 => "00110011",
 1718 => "01101011",
 1719 => "00100101",
 1720 => "10110111",
 1721 => "11110111",
 1722 => "01111010",
 1723 => "00101111",
 1724 => "10011011",
 1725 => "01111010",
 1726 => "00111001",
 1727 => "11101111",
 1728 => "01000110",
 1729 => "10100010",
 1730 => "10111011",
 1731 => "01001011",
 1732 => "10100110",
 1733 => "10101010",
 1734 => "10101011",
 1735 => "01000111",
 1736 => "01111000",
 1737 => "01111101",
 1738 => "01001011",
 1739 => "00010011",
 1740 => "10011011",
 1741 => "11010000",
 1742 => "11000010",
 1743 => "00011100",
 1744 => "01111100",
 1745 => "11011110",
 1746 => "01111001",
 1747 => "00100111",
 1748 => "00111011",
 1749 => "00111100",
 1750 => "01101101",
 1751 => "11001001",
 1752 => "10101111",
 1753 => "10101101",
 1754 => "11000110",
 1755 => "10101010",
 1756 => "00000010",
 1757 => "01001010",
 1758 => "01010001",
 1759 => "00101111",
 1760 => "00101001",
 1761 => "01000100",
 1762 => "11011101",
 1763 => "01101010",
 1764 => "10111100",
 1765 => "00001110",
 1766 => "01101100",
 1767 => "01101011",
 1768 => "11110011",
 1769 => "00100111",
 1770 => "11011001",
 1771 => "10001101",
 1772 => "00111100",
 1773 => "00001100",
 1774 => "11111010",
 1775 => "01010000",
 1776 => "11010101",
 1777 => "00011001",
 1778 => "01111011",
 1779 => "00010111",
 1780 => "01011111",
 1781 => "11000001",
 1782 => "10001101",
 1783 => "01000111",
 1784 => "00001110",
 1785 => "00010010",
 1786 => "11010000",
 1787 => "11111000",
 1788 => "01110110",
 1789 => "01010001",
 1790 => "01011111",
 1791 => "10111111",
 1792 => "01111001",
 1793 => "00001101",
 1794 => "11010101",
 1795 => "10000000",
 1796 => "00001010",
 1797 => "10110001",
 1798 => "11000111",
 1799 => "01001010",
 1800 => "01111100",
 1801 => "11100100",
 1802 => "11101100",
 1803 => "00111111",
 1804 => "00111100",
 1805 => "00101010",
 1806 => "11001011",
 1807 => "10100000",
 1808 => "01001110",
 1809 => "10100111",
 1810 => "10010000",
 1811 => "10010110",
 1812 => "01011000",
 1813 => "11010110",
 1814 => "00011100",
 1815 => "01111010",
 1816 => "10011001",
 1817 => "10000101",
 1818 => "10011001",
 1819 => "01000000",
 1820 => "10110011",
 1821 => "00000010",
 1822 => "01011001",
 1823 => "10110000",
 1824 => "01000101",
 1825 => "10000010",
 1826 => "11000001",
 1827 => "10110110",
 1828 => "00000000",
 1829 => "01100011",
 1830 => "01011110",
 1831 => "00001011",
 1832 => "00001101",
 1833 => "01000010",
 1834 => "00110100",
 1835 => "10000110",
 1836 => "10101010",
 1837 => "11000100",
 1838 => "11111001",
 1839 => "00011010",
 1840 => "11101010",
 1841 => "11101010",
 1842 => "01000101",
 1843 => "00000000",
 1844 => "00111001",
 1845 => "11100010",
 1846 => "11011100",
 1847 => "00001101",
 1848 => "11001110",
 1849 => "00111111",
 1850 => "00110011",
 1851 => "01101001",
 1852 => "10100101",
 1853 => "10101111",
 1854 => "00110111",
 1855 => "01101011",
 1856 => "11000101",
 1857 => "00111111",
 1858 => "11110111",
 1859 => "11000011",
 1860 => "10010010",
 1861 => "11100000",
 1862 => "11001111",
 1863 => "11101001",
 1864 => "01101010",
 1865 => "01011111",
 1866 => "01001110",
 1867 => "01011010",
 1868 => "10000000",
 1869 => "10111010",
 1870 => "11010110",
 1871 => "01101110",
 1872 => "00001011",
 1873 => "01001110",
 1874 => "01100100",
 1875 => "00110110",
 1876 => "01110001",
 1877 => "10011111",
 1878 => "01000001",
 1879 => "10000000",
 1880 => "00000110",
 1881 => "11001100",
 1882 => "01011000",
 1883 => "10010100",
 1884 => "01010101",
 1885 => "00011001",
 1886 => "10011110",
 1887 => "01111000",
 1888 => "01011010",
 1889 => "01010011",
 1890 => "00001111",
 1891 => "00001001",
 1892 => "00000110",
 1893 => "10010001",
 1894 => "10011011",
 1895 => "01101100",
 1896 => "00000000",
 1897 => "11011011",
 1898 => "11101110",
 1899 => "11011110",
 1900 => "10100001",
 1901 => "01110001",
 1902 => "11110010",
 1903 => "00000111",
 1904 => "01101111",
 1905 => "11010101",
 1906 => "01100111",
 1907 => "01011110",
 1908 => "00111101",
 1909 => "01011100",
 1910 => "11001001",
 1911 => "11111000",
 1912 => "01111100",
 1913 => "11110011",
 1914 => "10110000",
 1915 => "10100110",
 1916 => "10100010",
 1917 => "11011101",
 1918 => "00010101",
 1919 => "11000010",
 1920 => "01010010",
 1921 => "11101110",
 1922 => "00000001",
 1923 => "10110000",
 1924 => "01000100",
 1925 => "00001011",
 1926 => "00100110",
 1927 => "11100010",
 1928 => "11100001",
 1929 => "10100100",
 1930 => "00010110",
 1931 => "10001101",
 1932 => "10001000",
 1933 => "11010011",
 1934 => "10101101",
 1935 => "01111110",
 1936 => "10101100",
 1937 => "01110000",
 1938 => "00001000",
 1939 => "11110101",
 1940 => "00110111",
 1941 => "10011111",
 1942 => "11101100",
 1943 => "10010100",
 1944 => "11100011",
 1945 => "00101011",
 1946 => "11101101",
 1947 => "01110010",
 1948 => "10111110",
 1949 => "10000110",
 1950 => "01000010",
 1951 => "00110111",
 1952 => "00010111",
 1953 => "01011111",
 1954 => "10011101",
 1955 => "00000001",
 1956 => "01010100",
 1957 => "10100010",
 1958 => "11110101",
 1959 => "10110101",
 1960 => "11010100",
 1961 => "11100001",
 1962 => "11111110",
 1963 => "01110011",
 1964 => "10101100",
 1965 => "01111001",
 1966 => "01011101",
 1967 => "11110100",
 1968 => "00010111",
 1969 => "11111001",
 1970 => "00000010",
 1971 => "10100011",
 1972 => "10111001",
 1973 => "10100001",
 1974 => "11011010",
 1975 => "10100011",
 1976 => "11000100",
 1977 => "10010000",
 1978 => "01010111",
 1979 => "11011010",
 1980 => "00111001",
 1981 => "00100001",
 1982 => "00010000",
 1983 => "11000101",
 1984 => "00111000",
 1985 => "10010111",
 1986 => "10111010",
 1987 => "01010000",
 1988 => "01010001",
 1989 => "00000011",
 1990 => "10011000",
 1991 => "11000110",
 1992 => "00111001",
 1993 => "01001010",
 1994 => "00011011",
 1995 => "10111001",
 1996 => "10001000",
 1997 => "10111010",
 1998 => "00110101",
 1999 => "11011010",
 2000 => "10110011",
 2001 => "01100010",
 2002 => "10010110",
 2003 => "00000111",
 2004 => "01110101",
 2005 => "00101101",
 2006 => "10010000",
 2007 => "01010000",
 2008 => "10001110",
 2009 => "10101110",
 2010 => "01100111",
 2011 => "11000000",
 2012 => "01010000",
 2013 => "11010001",
 2014 => "01000011",
 2015 => "01111101",
 2016 => "10100100",
 2017 => "00000110",
 2018 => "00001001",
 2019 => "10001011",
 2020 => "11111100",
 2021 => "10000110",
 2022 => "11011001",
 2023 => "10101010",
 2024 => "11111010",
 2025 => "10011010",
 2026 => "00101101",
 2027 => "11110101",
 2028 => "01010010",
 2029 => "10010100",
 2030 => "11010110",
 2031 => "10011100",
 2032 => "10001000",
 2033 => "00100110",
 2034 => "11001011",
 2035 => "01000011",
 2036 => "01110000",
 2037 => "00100111",
 2038 => "11111101",
 2039 => "11000111",
 2040 => "01011000",
 2041 => "01101100",
 2042 => "10101011",
 2043 => "10101111",
 2044 => "10010010",
 2045 => "10100011",
 2046 => "00101010",
 2047 => "11001000",
 2048 => "10000101",
 2049 => "10011101",
 2050 => "01011001",
 2051 => "00010110",
 2052 => "00001111",
 2053 => "01001001",
 2054 => "11101001",
 2055 => "11100111",
 2056 => "01111101",
 2057 => "01100101",
 2058 => "01101111",
 2059 => "10001110",
 2060 => "10000001",
 2061 => "10110001",
 2062 => "00111001",
 2063 => "11100001",
 2064 => "00101000",
 2065 => "10111101",
 2066 => "00110111",
 2067 => "00100101",
 2068 => "10001001",
 2069 => "11100100",
 2070 => "01110110",
 2071 => "11100000",
 2072 => "10001110",
 2073 => "10111001",
 2074 => "01010010",
 2075 => "01010001",
 2076 => "10110010",
 2077 => "11001001",
 2078 => "10000110",
 2079 => "00010101",
 2080 => "11001100",
 2081 => "11010110",
 2082 => "01011100",
 2083 => "10100001",
 2084 => "11011100",
 2085 => "00011101",
 2086 => "01111000",
 2087 => "01101010",
 2088 => "00010100",
 2089 => "11011111",
 2090 => "01101001",
 2091 => "10011110",
 2092 => "00011110",
 2093 => "00000111",
 2094 => "01000100",
 2095 => "01000111",
 2096 => "00100010",
 2097 => "10011001",
 2098 => "11001100",
 2099 => "00000100",
 2100 => "01111110",
 2101 => "01001000",
 2102 => "00101101",
 2103 => "00011111",
 2104 => "01000110",
 2105 => "10010101",
 2106 => "11000111",
 2107 => "10000110",
 2108 => "10110001",
 2109 => "10010001",
 2110 => "10010101",
 2111 => "01010000",
 2112 => "11111101",
 2113 => "11011010",
 2114 => "10110111",
 2115 => "01110001",
 2116 => "11011110",
 2117 => "11000100",
 2118 => "00110010",
 2119 => "00111100",
 2120 => "01001001",
 2121 => "00100111",
 2122 => "00111001",
 2123 => "01011100",
 2124 => "00101000",
 2125 => "01000011",
 2126 => "11010011",
 2127 => "10110000",
 2128 => "00000111",
 2129 => "11111100",
 2130 => "01000111",
 2131 => "00011110",
 2132 => "01010001",
 2133 => "01011010",
 2134 => "00000010",
 2135 => "01110111",
 2136 => "10111000",
 2137 => "11100011",
 2138 => "00000011",
 2139 => "11000011",
 2140 => "11100001",
 2141 => "10001100",
 2142 => "00001010",
 2143 => "10010010",
 2144 => "00000011",
 2145 => "01100010",
 2146 => "10001110",
 2147 => "01111011",
 2148 => "10100111",
 2149 => "01100011",
 2150 => "01111001",
 2151 => "01100001",
 2152 => "10001000",
 2153 => "10100101",
 2154 => "01111100",
 2155 => "01011101",
 2156 => "11011011",
 2157 => "10111101",
 2158 => "00110011",
 2159 => "10111011",
 2160 => "00001111",
 2161 => "01111000",
 2162 => "10100100",
 2163 => "11100011",
 2164 => "10111010",
 2165 => "10100010",
 2166 => "11111101",
 2167 => "10011100",
 2168 => "11111110",
 2169 => "00101111",
 2170 => "11001000",
 2171 => "00111101",
 2172 => "11110010",
 2173 => "00101000",
 2174 => "00011111",
 2175 => "00101110",
 2176 => "00101000",
 2177 => "11110110",
 2178 => "00100111",
 2179 => "00010111",
 2180 => "10111000",
 2181 => "01110101",
 2182 => "10000101",
 2183 => "11001100",
 2184 => "10010101",
 2185 => "11011001",
 2186 => "01010101",
 2187 => "01011100",
 2188 => "10010011",
 2189 => "11010110",
 2190 => "01000001",
 2191 => "01111011",
 2192 => "10011001",
 2193 => "00001010",
 2194 => "00001000",
 2195 => "10110011",
 2196 => "01010001",
 2197 => "10100100",
 2198 => "10101010",
 2199 => "00111101",
 2200 => "10100010",
 2201 => "01000100",
 2202 => "01100110",
 2203 => "11100110",
 2204 => "00000000",
 2205 => "11011001",
 2206 => "00001010",
 2207 => "00101010",
 2208 => "00111101",
 2209 => "01110100",
 2210 => "00100000",
 2211 => "00110101",
 2212 => "01101110",
 2213 => "10111010",
 2214 => "00111001",
 2215 => "10000110",
 2216 => "00100010",
 2217 => "01101001",
 2218 => "10011110",
 2219 => "10000100",
 2220 => "10011001",
 2221 => "10110000",
 2222 => "10011110",
 2223 => "10111000",
 2224 => "01101011",
 2225 => "01111011",
 2226 => "11100001",
 2227 => "00101011",
 2228 => "10011100",
 2229 => "10101001",
 2230 => "10011110",
 2231 => "00101110",
 2232 => "11111110",
 2233 => "01011101",
 2234 => "10000111",
 2235 => "10011001",
 2236 => "00100011",
 2237 => "11001110",
 2238 => "10010100",
 2239 => "00100101",
 2240 => "00000101",
 2241 => "00110101",
 2242 => "10100100",
 2243 => "00100101",
 2244 => "11001110",
 2245 => "01000001",
 2246 => "10110110",
 2247 => "10100110",
 2248 => "11000110",
 2249 => "01111101",
 2250 => "00000100",
 2251 => "01101001",
 2252 => "11100101",
 2253 => "10110011",
 2254 => "10110101",
 2255 => "00110101",
 2256 => "11101010",
 2257 => "00000110",
 2258 => "00010001",
 2259 => "00011111",
 2260 => "01111010",
 2261 => "11111001",
 2262 => "11111011",
 2263 => "10001111",
 2264 => "11100100",
 2265 => "11000110",
 2266 => "10100010",
 2267 => "00110011",
 2268 => "11001101",
 2269 => "01101101",
 2270 => "01111000",
 2271 => "00101101",
 2272 => "10101001",
 2273 => "11110010",
 2274 => "10110010",
 2275 => "11111011",
 2276 => "01101000",
 2277 => "01110010",
 2278 => "10011000",
 2279 => "10110111",
 2280 => "10101011",
 2281 => "00111111",
 2282 => "10101101",
 2283 => "11001100",
 2284 => "01101101",
 2285 => "11100101",
 2286 => "11001000",
 2287 => "01010010",
 2288 => "11010101",
 2289 => "10100000",
 2290 => "11100100",
 2291 => "01011100",
 2292 => "00010011",
 2293 => "10010111",
 2294 => "01100010",
 2295 => "11000010",
 2296 => "00011100",
 2297 => "11010110",
 2298 => "10011011",
 2299 => "00100011",
 2300 => "11001011",
 2301 => "00001000",
 2302 => "10100001",
 2303 => "00010010",
 2304 => "01101001",
 2305 => "11111100",
 2306 => "00100110",
 2307 => "00010100",
 2308 => "11111000",
 2309 => "00000011",
 2310 => "00101000",
 2311 => "11001101",
 2312 => "01011101",
 2313 => "00111100",
 2314 => "00000100",
 2315 => "01110011",
 2316 => "00110000",
 2317 => "01111111",
 2318 => "11110000",
 2319 => "01110101",
 2320 => "10101111",
 2321 => "11011001",
 2322 => "00100101",
 2323 => "00101110",
 2324 => "11110011",
 2325 => "00010110",
 2326 => "01010110",
 2327 => "00100111",
 2328 => "00100001",
 2329 => "10101101",
 2330 => "00001010",
 2331 => "01100010",
 2332 => "00010100",
 2333 => "01011110",
 2334 => "11110011",
 2335 => "00000111",
 2336 => "11100001",
 2337 => "00100000",
 2338 => "10100010",
 2339 => "00010000",
 2340 => "00110011",
 2341 => "00111111",
 2342 => "11101001",
 2343 => "01101100",
 2344 => "00100011",
 2345 => "01110100",
 2346 => "11110110",
 2347 => "00101011",
 2348 => "00110011",
 2349 => "01111011",
 2350 => "11100000",
 2351 => "00010010",
 2352 => "10001010",
 2353 => "01110010",
 2354 => "10110111",
 2355 => "11001000",
 2356 => "00100001",
 2357 => "11000110",
 2358 => "01010000",
 2359 => "11001100",
 2360 => "10111100",
 2361 => "00111001",
 2362 => "00100010",
 2363 => "11010101",
 2364 => "00110010",
 2365 => "00001110",
 2366 => "11000000",
 2367 => "01100100",
 2368 => "01110010",
 2369 => "00010101",
 2370 => "11101101",
 2371 => "00010111",
 2372 => "01111011",
 2373 => "00101111",
 2374 => "01101011",
 2375 => "01001100",
 2376 => "11101101",
 2377 => "10011110",
 2378 => "01000100",
 2379 => "11111111",
 2380 => "01111110",
 2381 => "11110101",
 2382 => "00100001",
 2383 => "10011100",
 2384 => "11110001",
 2385 => "10001111",
 2386 => "11110100",
 2387 => "11111110",
 2388 => "11111001",
 2389 => "11000001",
 2390 => "11110101",
 2391 => "11001101",
 2392 => "00011001",
 2393 => "10111100",
 2394 => "01101110",
 2395 => "01010111",
 2396 => "10000100",
 2397 => "00000110",
 2398 => "11001111",
 2399 => "01101100",
 2400 => "01110001",
 2401 => "10011010",
 2402 => "11001101",
 2403 => "10110100",
 2404 => "00001100",
 2405 => "11011111",
 2406 => "10110110",
 2407 => "01111100",
 2408 => "11110110",
 2409 => "01110011",
 2410 => "10110110",
 2411 => "10001010",
 2412 => "10111001",
 2413 => "01011111",
 2414 => "10000001",
 2415 => "00001011",
 2416 => "10010100",
 2417 => "10010000",
 2418 => "10100101",
 2419 => "01101111",
 2420 => "11000111",
 2421 => "01010001",
 2422 => "00010001",
 2423 => "11000111",
 2424 => "01000111",
 2425 => "10000100",
 2426 => "01101111",
 2427 => "11111101",
 2428 => "01110000",
 2429 => "11000001",
 2430 => "01001001",
 2431 => "11111100",
 2432 => "01011101",
 2433 => "10011100",
 2434 => "11100010",
 2435 => "11100001",
 2436 => "01100101",
 2437 => "10101101",
 2438 => "11110111",
 2439 => "00110000",
 2440 => "00110100",
 2441 => "01001110",
 2442 => "01100110",
 2443 => "01011001",
 2444 => "11001000",
 2445 => "01101011",
 2446 => "11011001",
 2447 => "10011011",
 2448 => "00011011",
 2449 => "10000001",
 2450 => "01000000",
 2451 => "10111110",
 2452 => "11011011",
 2453 => "10101110",
 2454 => "10101010",
 2455 => "11100001",
 2456 => "01110110",
 2457 => "10000000",
 2458 => "10011101",
 2459 => "01101100",
 2460 => "00101111",
 2461 => "00111100",
 2462 => "01101111",
 2463 => "11001010",
 2464 => "10010100",
 2465 => "01000111",
 2466 => "01001110",
 2467 => "01000011",
 2468 => "10001011",
 2469 => "01111101",
 2470 => "01111101",
 2471 => "00101011",
 2472 => "01111010",
 2473 => "11000101",
 2474 => "01111001",
 2475 => "01101011",
 2476 => "10111100",
 2477 => "11100001",
 2478 => "11001001",
 2479 => "00011011",
 2480 => "11000110",
 2481 => "00111111",
 2482 => "10111111",
 2483 => "01001101",
 2484 => "00101001",
 2485 => "01010001",
 2486 => "00001011",
 2487 => "10001111",
 2488 => "01111000",
 2489 => "11100011",
 2490 => "01100110",
 2491 => "10101000",
 2492 => "00000101",
 2493 => "00000110",
 2494 => "01101100",
 2495 => "10101110",
 2496 => "10100001",
 2497 => "11110101",
 2498 => "11101011",
 2499 => "11000000",
 2500 => "11011110",
 2501 => "00110011",
 2502 => "01000100",
 2503 => "10110001",
 2504 => "10111011",
 2505 => "01110000",
 2506 => "00001011",
 2507 => "00101100",
 2508 => "00111001",
 2509 => "00111110",
 2510 => "11100111",
 2511 => "00100110",
 2512 => "11001110",
 2513 => "00011101",
 2514 => "11010100",
 2515 => "01010011",
 2516 => "11010010",
 2517 => "00000000",
 2518 => "00111110",
 2519 => "00011100",
 2520 => "01001010",
 2521 => "01010010",
 2522 => "10011001",
 2523 => "11110111",
 2524 => "00010110",
 2525 => "01100111",
 2526 => "00101001",
 2527 => "00011111",
 2528 => "00110110",
 2529 => "01100001",
 2530 => "01111000",
 2531 => "11011010",
 2532 => "11111100",
 2533 => "10111100",
 2534 => "10100111",
 2535 => "11101110",
 2536 => "11000101",
 2537 => "11111001",
 2538 => "00010101",
 2539 => "01001011",
 2540 => "10000110",
 2541 => "00011110",
 2542 => "00010011",
 2543 => "11111011",
 2544 => "01110100",
 2545 => "10001011",
 2546 => "11001110",
 2547 => "10100100",
 2548 => "00001011",
 2549 => "01011011",
 2550 => "00110001",
 2551 => "10000111",
 2552 => "01100010",
 2553 => "00101100",
 2554 => "10110110",
 2555 => "10111110",
 2556 => "00011001",
 2557 => "00010010",
 2558 => "00100000",
 2559 => "01011101",
 2560 => "11111000",
 2561 => "10101110",
 2562 => "01000100",
 2563 => "01011100",
 2564 => "01001010",
 2565 => "01011001",
 2566 => "01100011",
 2567 => "10011110",
 2568 => "10101101",
 2569 => "00011011",
 2570 => "11001010",
 2571 => "10101000",
 2572 => "11001000",
 2573 => "01101010",
 2574 => "11011100",
 2575 => "01011000",
 2576 => "00001010",
 2577 => "10111010",
 2578 => "00001000",
 2579 => "00111001",
 2580 => "10000000",
 2581 => "10011000",
 2582 => "11011101",
 2583 => "00100010",
 2584 => "00100101",
 2585 => "00010011",
 2586 => "00101111",
 2587 => "01101100",
 2588 => "01001010",
 2589 => "10100000",
 2590 => "11000101",
 2591 => "11001010",
 2592 => "01010000",
 2593 => "10000011",
 2594 => "10001010",
 2595 => "11110000",
 2596 => "00111100",
 2597 => "00011110",
 2598 => "00100001",
 2599 => "01001001",
 2600 => "11001110",
 2601 => "11101000",
 2602 => "10111010",
 2603 => "11001011",
 2604 => "01111010",
 2605 => "00001011",
 2606 => "00100110",
 2607 => "11111001",
 2608 => "11101011",
 2609 => "01101010",
 2610 => "10111100",
 2611 => "10010011",
 2612 => "10111100",
 2613 => "11110111",
 2614 => "11011101",
 2615 => "10110111",
 2616 => "11011110",
 2617 => "00011011",
 2618 => "00010000",
 2619 => "11110010",
 2620 => "01101010",
 2621 => "01110101",
 2622 => "10100010",
 2623 => "00111110",
 2624 => "10101110",
 2625 => "10010000",
 2626 => "01110011",
 2627 => "00101011",
 2628 => "00011101",
 2629 => "11000000",
 2630 => "11001010",
 2631 => "11000000",
 2632 => "11101001",
 2633 => "11001010",
 2634 => "10110000",
 2635 => "11010110",
 2636 => "11111101",
 2637 => "01010011",
 2638 => "00111000",
 2639 => "11101010",
 2640 => "00001000",
 2641 => "10010001",
 2642 => "10111101",
 2643 => "01100000",
 2644 => "10010110",
 2645 => "00100001",
 2646 => "00101000",
 2647 => "11111010",
 2648 => "10001100",
 2649 => "10010011",
 2650 => "00111101",
 2651 => "01101110",
 2652 => "11001001",
 2653 => "01001011",
 2654 => "11011011",
 2655 => "01111000",
 2656 => "10101011",
 2657 => "11010111",
 2658 => "10111100",
 2659 => "01010010",
 2660 => "10100000",
 2661 => "10001100",
 2662 => "11000011",
 2663 => "10101110",
 2664 => "00010111",
 2665 => "01000110",
 2666 => "11101101",
 2667 => "11000010",
 2668 => "01011000",
 2669 => "10110101",
 2670 => "11100100",
 2671 => "10001010",
 2672 => "10000010",
 2673 => "00001101",
 2674 => "10111100",
 2675 => "10001000",
 2676 => "11010001",
 2677 => "01001100",
 2678 => "11001011",
 2679 => "11000111",
 2680 => "00000001",
 2681 => "00000000",
 2682 => "11110011",
 2683 => "00010010",
 2684 => "01011000",
 2685 => "11111111",
 2686 => "00111010",
 2687 => "00110000",
 2688 => "00111001",
 2689 => "11000111",
 2690 => "00101000",
 2691 => "11001111",
 2692 => "01111111",
 2693 => "01000111",
 2694 => "00111011",
 2695 => "00011101",
 2696 => "11000111",
 2697 => "10110110",
 2698 => "00100011",
 2699 => "11111110",
 2700 => "10101100",
 2701 => "10010100",
 2702 => "01010100",
 2703 => "00011100",
 2704 => "00110011",
 2705 => "11110011",
 2706 => "11101111",
 2707 => "10111111",
 2708 => "11001000",
 2709 => "10111000",
 2710 => "00011011",
 2711 => "00101111",
 2712 => "11010010",
 2713 => "01101101",
 2714 => "00001010",
 2715 => "10101000",
 2716 => "00100101",
 2717 => "00101111",
 2718 => "01110001",
 2719 => "11001101",
 2720 => "01110000",
 2721 => "10001110",
 2722 => "00110101",
 2723 => "10011101",
 2724 => "00001100",
 2725 => "11110010",
 2726 => "10100100",
 2727 => "00010100",
 2728 => "00010010",
 2729 => "10011100",
 2730 => "11001111",
 2731 => "01110110",
 2732 => "01000011",
 2733 => "00110010",
 2734 => "00001100",
 2735 => "01010101",
 2736 => "00101101",
 2737 => "11111100",
 2738 => "01100000",
 2739 => "10001110",
 2740 => "11111000",
 2741 => "10010011",
 2742 => "01101000",
 2743 => "11011111",
 2744 => "11101000",
 2745 => "10101011",
 2746 => "11010001",
 2747 => "00001011",
 2748 => "10011100",
 2749 => "11001011",
 2750 => "00101000",
 2751 => "00110001",
 2752 => "11111010",
 2753 => "10100111",
 2754 => "11011001",
 2755 => "00000011",
 2756 => "10111011",
 2757 => "10111100",
 2758 => "00110100",
 2759 => "01010100",
 2760 => "11100111",
 2761 => "11011010",
 2762 => "00100101",
 2763 => "00010011",
 2764 => "00110010",
 2765 => "11111010",
 2766 => "00100111",
 2767 => "00011010",
 2768 => "11010101",
 2769 => "11000010",
 2770 => "01011111",
 2771 => "00001001",
 2772 => "01101101",
 2773 => "10110010",
 2774 => "11000000",
 2775 => "11101110",
 2776 => "00100100",
 2777 => "10111110",
 2778 => "01001101",
 2779 => "10111101",
 2780 => "10010101",
 2781 => "00010001",
 2782 => "10001011",
 2783 => "01011000",
 2784 => "00111110",
 2785 => "00100001",
 2786 => "01110100",
 2787 => "01100110",
 2788 => "00010100",
 2789 => "00011101",
 2790 => "01111101",
 2791 => "00100110",
 2792 => "11101010",
 2793 => "00101111",
 2794 => "11100000",
 2795 => "10010000",
 2796 => "11100000",
 2797 => "10100101",
 2798 => "01110010",
 2799 => "10100100",
 2800 => "01111001",
 2801 => "01101101",
 2802 => "10010110",
 2803 => "11110100",
 2804 => "10001100",
 2805 => "01110110",
 2806 => "01111011",
 2807 => "00100110",
 2808 => "11011011",
 2809 => "11000110",
 2810 => "11010101",
 2811 => "10010000",
 2812 => "00111011",
 2813 => "01101111",
 2814 => "11110101",
 2815 => "10110001",
 2816 => "01111011",
 2817 => "10100100",
 2818 => "11110111",
 2819 => "11101010",
 2820 => "01010101",
 2821 => "11010011",
 2822 => "00011000",
 2823 => "11110000",
 2824 => "11000101",
 2825 => "11010001",
 2826 => "11000001",
 2827 => "01110101",
 2828 => "01000011",
 2829 => "01010101",
 2830 => "00101001",
 2831 => "10011111",
 2832 => "11011100",
 2833 => "10110101",
 2834 => "11111110",
 2835 => "01110111",
 2836 => "11111100",
 2837 => "10000011",
 2838 => "11001010",
 2839 => "00010011",
 2840 => "00110000",
 2841 => "10101000",
 2842 => "01101110",
 2843 => "11101011",
 2844 => "11100010",
 2845 => "00100011",
 2846 => "11000111",
 2847 => "10101100",
 2848 => "00010101",
 2849 => "10101110",
 2850 => "01000001",
 2851 => "01100100",
 2852 => "01110100",
 2853 => "11100000",
 2854 => "01100010",
 2855 => "11000100",
 2856 => "00101110",
 2857 => "11001010",
 2858 => "11000001",
 2859 => "00101001",
 2860 => "11000111",
 2861 => "11100111",
 2862 => "00111000",
 2863 => "11100100",
 2864 => "11010110",
 2865 => "10111101",
 2866 => "01100111",
 2867 => "11011100",
 2868 => "01001011",
 2869 => "00011101",
 2870 => "11100001",
 2871 => "00110001",
 2872 => "00111011",
 2873 => "11000110",
 2874 => "10100110",
 2875 => "11110101",
 2876 => "00010001",
 2877 => "00101111",
 2878 => "11101001",
 2879 => "01100111",
 2880 => "01101101",
 2881 => "11000111",
 2882 => "00001101",
 2883 => "00001111",
 2884 => "10011000",
 2885 => "10101001",
 2886 => "01010001",
 2887 => "11110101",
 2888 => "11110111",
 2889 => "11100011",
 2890 => "01101110",
 2891 => "11100000",
 2892 => "11110001",
 2893 => "10100011",
 2894 => "10100110",
 2895 => "11001111",
 2896 => "01011011",
 2897 => "11001010",
 2898 => "10000111",
 2899 => "10101000",
 2900 => "01111101",
 2901 => "10111011",
 2902 => "11111111",
 2903 => "00010010",
 2904 => "00111001",
 2905 => "01000100",
 2906 => "10011011",
 2907 => "01111100",
 2908 => "00000010",
 2909 => "01110001",
 2910 => "00000111",
 2911 => "10101000",
 2912 => "10001010",
 2913 => "10000101",
 2914 => "00010000",
 2915 => "00101001",
 2916 => "00010010",
 2917 => "11011001",
 2918 => "11101001",
 2919 => "10100010",
 2920 => "11010101",
 2921 => "11001111",
 2922 => "01111001",
 2923 => "10001110",
 2924 => "00101111",
 2925 => "01101100",
 2926 => "10000000",
 2927 => "11000010",
 2928 => "11010100",
 2929 => "10011101",
 2930 => "10110111",
 2931 => "01100010",
 2932 => "11101110",
 2933 => "01000001",
 2934 => "00010110",
 2935 => "01001111",
 2936 => "10111010",
 2937 => "11010011",
 2938 => "10101001",
 2939 => "11110010",
 2940 => "01100000",
 2941 => "11010110",
 2942 => "10000111",
 2943 => "10111010",
 2944 => "11111010",
 2945 => "10100100",
 2946 => "00011010",
 2947 => "10001010",
 2948 => "10001110",
 2949 => "00010011",
 2950 => "11111110",
 2951 => "01001010",
 2952 => "10001101",
 2953 => "00000000",
 2954 => "11010011",
 2955 => "10000011",
 2956 => "10111110",
 2957 => "11111111",
 2958 => "11101001",
 2959 => "10011010",
 2960 => "00010110",
 2961 => "00000010",
 2962 => "11101100",
 2963 => "11011100",
 2964 => "00000111",
 2965 => "10100100",
 2966 => "10101000",
 2967 => "11101001",
 2968 => "10010100",
 2969 => "01001000",
 2970 => "01111000",
 2971 => "10111010",
 2972 => "11001111",
 2973 => "11110100",
 2974 => "01111110",
 2975 => "10001111",
 2976 => "00011000",
 2977 => "01001100",
 2978 => "01010100",
 2979 => "01110001",
 2980 => "01010100",
 2981 => "11111001",
 2982 => "01000010",
 2983 => "10001010",
 2984 => "10110001",
 2985 => "11111100",
 2986 => "00111100",
 2987 => "11001000",
 2988 => "11001101",
 2989 => "10000110",
 2990 => "11001111",
 2991 => "10101010",
 2992 => "01011000",
 2993 => "00010000",
 2994 => "01110101",
 2995 => "10010011",
 2996 => "00111011",
 2997 => "01100011",
 2998 => "00111001",
 2999 => "01001001",
 3000 => "10100010",
 3001 => "00011111",
 3002 => "01001100",
 3003 => "10111101",
 3004 => "11101011",
 3005 => "11111101",
 3006 => "00111111",
 3007 => "00110100",
 3008 => "01101100",
 3009 => "11001101",
 3010 => "01110100",
 3011 => "11110110",
 3012 => "00001110",
 3013 => "01010101",
 3014 => "10001111",
 3015 => "01111010",
 3016 => "01111001",
 3017 => "11101010",
 3018 => "10110011",
 3019 => "10110101",
 3020 => "00101101",
 3021 => "10000111",
 3022 => "00110000",
 3023 => "00111110",
 3024 => "00000101",
 3025 => "11100100",
 3026 => "10000010",
 3027 => "10110001",
 3028 => "11001011",
 3029 => "10111000",
 3030 => "00111010",
 3031 => "00100000",
 3032 => "01011100",
 3033 => "00101000",
 3034 => "00001000",
 3035 => "10111010",
 3036 => "01111010",
 3037 => "01000011",
 3038 => "00000110",
 3039 => "00111000",
 3040 => "11011001",
 3041 => "10000001",
 3042 => "01001110",
 3043 => "11001100",
 3044 => "11010010",
 3045 => "10001010",
 3046 => "01011101",
 3047 => "11001000",
 3048 => "00011101",
 3049 => "00101101",
 3050 => "10100111",
 3051 => "00111000",
 3052 => "01010011",
 3053 => "00101100",
 3054 => "00111011",
 3055 => "11110010",
 3056 => "11111111",
 3057 => "11110100",
 3058 => "10101000",
 3059 => "10101010",
 3060 => "10011011",
 3061 => "00101001",
 3062 => "11010010",
 3063 => "11111111",
 3064 => "10010111",
 3065 => "01101100",
 3066 => "11001011",
 3067 => "01110110",
 3068 => "00111111",
 3069 => "10110000",
 3070 => "00100011",
 3071 => "11001110",
 3072 => "11000000",
 3073 => "10110100",
 3074 => "00011001",
 3075 => "10001011",
 3076 => "10111110",
 3077 => "01110011",
 3078 => "01110101",
 3079 => "00001000",
 3080 => "11000100",
 3081 => "00100001",
 3082 => "10000100",
 3083 => "00111011",
 3084 => "00110000",
 3085 => "11110110",
 3086 => "00010000",
 3087 => "11001000",
 3088 => "00001101",
 3089 => "11000000",
 3090 => "11001001",
 3091 => "00110100",
 3092 => "10010011",
 3093 => "00001010",
 3094 => "11000011",
 3095 => "10001100",
 3096 => "00010010",
 3097 => "11101010",
 3098 => "00111010",
 3099 => "10000001",
 3100 => "11110111",
 3101 => "11111000",
 3102 => "10111000",
 3103 => "11101010",
 3104 => "10100000",
 3105 => "11101101",
 3106 => "01100010",
 3107 => "00001001",
 3108 => "00011111",
 3109 => "01000111",
 3110 => "00110110",
 3111 => "10000010",
 3112 => "11101111",
 3113 => "10110010",
 3114 => "11011100",
 3115 => "00000101",
 3116 => "01100010",
 3117 => "11110011",
 3118 => "00011010",
 3119 => "10011011",
 3120 => "01100000",
 3121 => "11100101",
 3122 => "01101010",
 3123 => "00000110",
 3124 => "11100110",
 3125 => "11001010",
 3126 => "01111010",
 3127 => "11110010",
 3128 => "01101101",
 3129 => "10011011",
 3130 => "10111100",
 3131 => "10110000",
 3132 => "00111101",
 3133 => "11101010",
 3134 => "00010101",
 3135 => "00010111",
 3136 => "01011100",
 3137 => "00111101",
 3138 => "11000111",
 3139 => "01010000",
 3140 => "01011110",
 3141 => "10100100",
 3142 => "10100011",
 3143 => "00000101",
 3144 => "11100011",
 3145 => "00011011",
 3146 => "00101101",
 3147 => "10000010",
 3148 => "10010100",
 3149 => "11111011",
 3150 => "01010001",
 3151 => "10011010",
 3152 => "11101001",
 3153 => "10010001",
 3154 => "10101101",
 3155 => "11011100",
 3156 => "10011100",
 3157 => "01000110",
 3158 => "01111100",
 3159 => "11010110",
 3160 => "10101010",
 3161 => "01000010",
 3162 => "10011100",
 3163 => "01001110",
 3164 => "10011011",
 3165 => "11000000",
 3166 => "11111101",
 3167 => "10000011",
 3168 => "00000010",
 3169 => "11001110",
 3170 => "00110000",
 3171 => "10001000",
 3172 => "11011000",
 3173 => "01011100",
 3174 => "00010000",
 3175 => "01110101",
 3176 => "00100010",
 3177 => "01110100",
 3178 => "11111000",
 3179 => "01011011",
 3180 => "01011110",
 3181 => "10010111",
 3182 => "01111001",
 3183 => "10000010",
 3184 => "01101100",
 3185 => "01101010",
 3186 => "00010110",
 3187 => "00011011",
 3188 => "10101011",
 3189 => "01001110",
 3190 => "01100111",
 3191 => "01011111",
 3192 => "10101010",
 3193 => "10010110",
 3194 => "11011001",
 3195 => "10000000",
 3196 => "00100110",
 3197 => "10110011",
 3198 => "11000011",
 3199 => "00000010",
 3200 => "11111110",
 3201 => "11110011",
 3202 => "10001011",
 3203 => "11101110",
 3204 => "00101001",
 3205 => "11111010",
 3206 => "10010001",
 3207 => "01000011",
 3208 => "11011111",
 3209 => "10011001",
 3210 => "00101000",
 3211 => "11011110",
 3212 => "11001000",
 3213 => "11101011",
 3214 => "10011110",
 3215 => "01110000",
 3216 => "10000101",
 3217 => "10100110",
 3218 => "00011010",
 3219 => "00100101",
 3220 => "00111011",
 3221 => "10000110",
 3222 => "11001111",
 3223 => "01001110",
 3224 => "11011011",
 3225 => "01011100",
 3226 => "10010000",
 3227 => "10001110",
 3228 => "00011111",
 3229 => "11101101",
 3230 => "01011100",
 3231 => "01011011",
 3232 => "11010000",
 3233 => "11000001",
 3234 => "01011000",
 3235 => "00100110",
 3236 => "01010111",
 3237 => "10010110",
 3238 => "00110110",
 3239 => "10110000",
 3240 => "01110010",
 3241 => "10111010",
 3242 => "11101000",
 3243 => "01001110",
 3244 => "01010011",
 3245 => "11100000",
 3246 => "11110100",
 3247 => "10100000",
 3248 => "11011110",
 3249 => "11100010",
 3250 => "11010000",
 3251 => "11111100",
 3252 => "10000011",
 3253 => "00111111",
 3254 => "11001010",
 3255 => "00100011",
 3256 => "01000100",
 3257 => "10010000",
 3258 => "01111001",
 3259 => "11100001",
 3260 => "00001100",
 3261 => "01000010",
 3262 => "01111110",
 3263 => "10111101",
 3264 => "11111101",
 3265 => "11010010",
 3266 => "00000010",
 3267 => "11000101",
 3268 => "10011111",
 3269 => "00100011",
 3270 => "11000110",
 3271 => "00010011",
 3272 => "10101111",
 3273 => "01100111",
 3274 => "10100001",
 3275 => "00111101",
 3276 => "01110010",
 3277 => "11111111",
 3278 => "00110100",
 3279 => "10010010",
 3280 => "00001010",
 3281 => "01011000",
 3282 => "01101111",
 3283 => "00001011",
 3284 => "11111101",
 3285 => "01001010",
 3286 => "11111111",
 3287 => "10110110",
 3288 => "10110100",
 3289 => "00110100",
 3290 => "11000101",
 3291 => "10000000",
 3292 => "11101011",
 3293 => "00010111",
 3294 => "10001000",
 3295 => "00000011",
 3296 => "01111001",
 3297 => "00010110",
 3298 => "00110110",
 3299 => "01101100",
 3300 => "01110000",
 3301 => "10000000",
 3302 => "10001101",
 3303 => "00011010",
 3304 => "11011011",
 3305 => "00010000",
 3306 => "00001100",
 3307 => "00001110",
 3308 => "11001000",
 3309 => "11100010",
 3310 => "11010000",
 3311 => "00111000",
 3312 => "00011101",
 3313 => "11100111",
 3314 => "10000011",
 3315 => "00110001",
 3316 => "11110111",
 3317 => "00100001",
 3318 => "01011011",
 3319 => "11010111",
 3320 => "01010111",
 3321 => "00100001",
 3322 => "01001011",
 3323 => "10000110",
 3324 => "10101110",
 3325 => "10010010",
 3326 => "01111110",
 3327 => "10011111",
 3328 => "00011100",
 3329 => "11100101",
 3330 => "01110011",
 3331 => "10110001",
 3332 => "11100010",
 3333 => "01001011",
 3334 => "01101011",
 3335 => "01111100",
 3336 => "01110000",
 3337 => "11110110",
 3338 => "11011010",
 3339 => "11011000",
 3340 => "00010100",
 3341 => "01111100",
 3342 => "11110001",
 3343 => "11101101",
 3344 => "10111000",
 3345 => "11110100",
 3346 => "01111111",
 3347 => "10010100",
 3348 => "00101111",
 3349 => "01001001",
 3350 => "11000000",
 3351 => "11101010",
 3352 => "00011111",
 3353 => "11000001",
 3354 => "00100011",
 3355 => "01000100",
 3356 => "01110110",
 3357 => "00001101",
 3358 => "00110000",
 3359 => "01110100",
 3360 => "10011010",
 3361 => "11011110",
 3362 => "11100011",
 3363 => "00000010",
 3364 => "10100110",
 3365 => "11011000",
 3366 => "01111110",
 3367 => "00000001",
 3368 => "11011000",
 3369 => "11111001",
 3370 => "11000110",
 3371 => "10101111",
 3372 => "11010101",
 3373 => "00010111",
 3374 => "00001100",
 3375 => "01111010",
 3376 => "11100011",
 3377 => "01110010",
 3378 => "00100111",
 3379 => "00110011",
 3380 => "11110100",
 3381 => "11011111",
 3382 => "00110110",
 3383 => "00110010",
 3384 => "00001010",
 3385 => "11110001",
 3386 => "01011110",
 3387 => "10111010",
 3388 => "01110000",
 3389 => "01110110",
 3390 => "10011011",
 3391 => "10001001",
 3392 => "10011110",
 3393 => "00111000",
 3394 => "10110100",
 3395 => "10001001",
 3396 => "00100010",
 3397 => "01111010",
 3398 => "01011111",
 3399 => "00001111",
 3400 => "01111110",
 3401 => "11001101",
 3402 => "11010001",
 3403 => "10010111",
 3404 => "01010100",
 3405 => "10111011",
 3406 => "01110100",
 3407 => "00000001",
 3408 => "01010101",
 3409 => "11001010",
 3410 => "01000100",
 3411 => "01100000",
 3412 => "11101010",
 3413 => "01100001",
 3414 => "00000101",
 3415 => "11111011",
 3416 => "01110101",
 3417 => "11000011",
 3418 => "01000101",
 3419 => "01010111",
 3420 => "10100001",
 3421 => "10100001",
 3422 => "11110011",
 3423 => "10110010",
 3424 => "11100011",
 3425 => "11101100",
 3426 => "11101000",
 3427 => "00010100",
 3428 => "01001100",
 3429 => "10011011",
 3430 => "11000111",
 3431 => "11001110",
 3432 => "10100010",
 3433 => "10111001",
 3434 => "01001111",
 3435 => "00111001",
 3436 => "00001010",
 3437 => "01111010",
 3438 => "01100011",
 3439 => "10011100",
 3440 => "11110101",
 3441 => "11001111",
 3442 => "11111111",
 3443 => "00110101",
 3444 => "00110000",
 3445 => "01111111",
 3446 => "00100000",
 3447 => "10000100",
 3448 => "11100001",
 3449 => "10110111",
 3450 => "11110011",
 3451 => "00100100",
 3452 => "01110110",
 3453 => "10110000",
 3454 => "11000000",
 3455 => "11000011",
 3456 => "01001001",
 3457 => "00110110",
 3458 => "00001000",
 3459 => "11000010",
 3460 => "10001000",
 3461 => "01111101",
 3462 => "01111111",
 3463 => "10011110",
 3464 => "11001000",
 3465 => "11001000",
 3466 => "11010001",
 3467 => "01110011",
 3468 => "00001000",
 3469 => "11010100",
 3470 => "00111100",
 3471 => "11110111",
 3472 => "01010100",
 3473 => "11101000",
 3474 => "11000011",
 3475 => "11010000",
 3476 => "11001111",
 3477 => "11001101",
 3478 => "00000111",
 3479 => "00111110",
 3480 => "00100101",
 3481 => "01101000",
 3482 => "10010101",
 3483 => "10010011",
 3484 => "00001101",
 3485 => "10011111",
 3486 => "11100100",
 3487 => "10101001",
 3488 => "11010001",
 3489 => "11110010",
 3490 => "00100001",
 3491 => "00000001",
 3492 => "11110111",
 3493 => "10001110",
 3494 => "11001000",
 3495 => "11000011",
 3496 => "10100111",
 3497 => "11010000",
 3498 => "10110111",
 3499 => "00100111",
 3500 => "10011101",
 3501 => "10100011",
 3502 => "00011110",
 3503 => "01100111",
 3504 => "00010010",
 3505 => "10101010",
 3506 => "00000000",
 3507 => "00011100",
 3508 => "11010000",
 3509 => "01110010",
 3510 => "10110101",
 3511 => "11100000",
 3512 => "01000100",
 3513 => "01010101",
 3514 => "11111110",
 3515 => "01111101",
 3516 => "01010100",
 3517 => "00011001",
 3518 => "01010111",
 3519 => "01101001",
 3520 => "01010111",
 3521 => "00101100",
 3522 => "01101111",
 3523 => "01000001",
 3524 => "00001110",
 3525 => "01101000",
 3526 => "01010101",
 3527 => "01110111",
 3528 => "00000111",
 3529 => "11100110",
 3530 => "01110011",
 3531 => "00110010",
 3532 => "00001110",
 3533 => "01100011",
 3534 => "00100000",
 3535 => "11011011",
 3536 => "01010101",
 3537 => "01101101",
 3538 => "10010110",
 3539 => "10101100",
 3540 => "00100011",
 3541 => "00010100",
 3542 => "00111011",
 3543 => "10110001",
 3544 => "10100001",
 3545 => "01110101",
 3546 => "00110011",
 3547 => "10001010",
 3548 => "01101100",
 3549 => "01100111",
 3550 => "10100101",
 3551 => "10011011",
 3552 => "11010101",
 3553 => "10111101",
 3554 => "00010011",
 3555 => "10110100",
 3556 => "10101111",
 3557 => "10001001",
 3558 => "11011010",
 3559 => "01010100",
 3560 => "00011001",
 3561 => "10000111",
 3562 => "10000011",
 3563 => "00000100",
 3564 => "00111110",
 3565 => "01101000",
 3566 => "00100110",
 3567 => "00010011",
 3568 => "01110001",
 3569 => "10010001",
 3570 => "11011001",
 3571 => "01111000",
 3572 => "11110110",
 3573 => "01111000",
 3574 => "10100101",
 3575 => "10100011",
 3576 => "10011100",
 3577 => "11101101",
 3578 => "00011001",
 3579 => "00010111",
 3580 => "00010110",
 3581 => "00000101",
 3582 => "11001101",
 3583 => "11010100",
 3584 => "10011001",
 3585 => "11111001",
 3586 => "10111100",
 3587 => "01111111",
 3588 => "11100010",
 3589 => "11011111",
 3590 => "00101101",
 3591 => "11111111",
 3592 => "01011000",
 3593 => "10011100",
 3594 => "10000001",
 3595 => "11111100",
 3596 => "10101010",
 3597 => "00100010",
 3598 => "00110111",
 3599 => "11000100",
 3600 => "10100100",
 3601 => "10001101",
 3602 => "11111101",
 3603 => "00100110",
 3604 => "01110001",
 3605 => "00000011",
 3606 => "10010101",
 3607 => "00100100",
 3608 => "01000010",
 3609 => "10101110",
 3610 => "10011001",
 3611 => "01100100",
 3612 => "01110000",
 3613 => "00110001",
 3614 => "10001100",
 3615 => "11100101",
 3616 => "10001010",
 3617 => "10001101",
 3618 => "11111100",
 3619 => "11100100",
 3620 => "11110010",
 3621 => "10000001",
 3622 => "11010101",
 3623 => "10100001",
 3624 => "10000111",
 3625 => "11001100",
 3626 => "00000010",
 3627 => "10111011",
 3628 => "00101011",
 3629 => "11101000",
 3630 => "00101000",
 3631 => "10010001",
 3632 => "00001110",
 3633 => "01000110",
 3634 => "10111011",
 3635 => "11101010",
 3636 => "00110100",
 3637 => "11111111",
 3638 => "10100101",
 3639 => "00011010",
 3640 => "10010010",
 3641 => "00101010",
 3642 => "00111000",
 3643 => "00000000",
 3644 => "11000000",
 3645 => "00100101",
 3646 => "01000100",
 3647 => "00101011",
 3648 => "10110000",
 3649 => "00100110",
 3650 => "01011001",
 3651 => "11111000",
 3652 => "00100000",
 3653 => "01000010",
 3654 => "01100101",
 3655 => "01011001",
 3656 => "11000001",
 3657 => "01100101",
 3658 => "00101001",
 3659 => "10111000",
 3660 => "00110011",
 3661 => "10101111",
 3662 => "11011101",
 3663 => "00110110",
 3664 => "11110100",
 3665 => "01111001",
 3666 => "11111110",
 3667 => "01100110",
 3668 => "01110000",
 3669 => "00000001",
 3670 => "00001010",
 3671 => "10110010",
 3672 => "10100010",
 3673 => "11010001",
 3674 => "00001001",
 3675 => "10011100",
 3676 => "11110001",
 3677 => "00001101",
 3678 => "10001101",
 3679 => "00010011",
 3680 => "00001001",
 3681 => "11110011",
 3682 => "11110000",
 3683 => "00100000",
 3684 => "10100111",
 3685 => "11000100",
 3686 => "11001101",
 3687 => "00100001",
 3688 => "00111000",
 3689 => "11110010",
 3690 => "11011110",
 3691 => "11011111",
 3692 => "01011010",
 3693 => "00110000",
 3694 => "11000100",
 3695 => "10111101",
 3696 => "00100011",
 3697 => "10000100",
 3698 => "01100011",
 3699 => "00010000",
 3700 => "10101110",
 3701 => "01100001",
 3702 => "11100011",
 3703 => "01001100",
 3704 => "10110100",
 3705 => "11000010",
 3706 => "01011011",
 3707 => "01010111",
 3708 => "10100100",
 3709 => "11101011",
 3710 => "00111001",
 3711 => "10101111",
 3712 => "11011001",
 3713 => "11101111",
 3714 => "00011010",
 3715 => "01100111",
 3716 => "10010010",
 3717 => "01110100",
 3718 => "10111111",
 3719 => "10100010",
 3720 => "01001010",
 3721 => "10110110",
 3722 => "01001111",
 3723 => "11100000",
 3724 => "01011001",
 3725 => "01000110",
 3726 => "00011111",
 3727 => "01110111",
 3728 => "01001100",
 3729 => "00001001",
 3730 => "01000010",
 3731 => "01110110",
 3732 => "10100111",
 3733 => "11000110",
 3734 => "10110101",
 3735 => "00010001",
 3736 => "00001011",
 3737 => "00000111",
 3738 => "01111010",
 3739 => "10100101",
 3740 => "11111110",
 3741 => "11111110",
 3742 => "00110001",
 3743 => "01010101",
 3744 => "01011010",
 3745 => "01110110",
 3746 => "01001110",
 3747 => "01000111",
 3748 => "00110010",
 3749 => "01110101",
 3750 => "11100100",
 3751 => "01100111",
 3752 => "00001011",
 3753 => "00100100",
 3754 => "10000111",
 3755 => "10000010",
 3756 => "00110100",
 3757 => "00100100",
 3758 => "01011011",
 3759 => "11010101",
 3760 => "10001111",
 3761 => "10011111",
 3762 => "10001001",
 3763 => "11100100",
 3764 => "00011101",
 3765 => "00110111",
 3766 => "10001010",
 3767 => "00100100",
 3768 => "01111001",
 3769 => "10001100",
 3770 => "10011010",
 3771 => "11001001",
 3772 => "10101101",
 3773 => "00000110",
 3774 => "10101101",
 3775 => "10010110",
 3776 => "01110111",
 3777 => "00000100",
 3778 => "00111001",
 3779 => "00110110",
 3780 => "01111110",
 3781 => "11000010",
 3782 => "10101100",
 3783 => "01110001",
 3784 => "10010100",
 3785 => "10110100",
 3786 => "11011011",
 3787 => "10100010",
 3788 => "10101010",
 3789 => "10111110",
 3790 => "10110100",
 3791 => "10011010",
 3792 => "00011011",
 3793 => "11110001",
 3794 => "00001010",
 3795 => "01101011",
 3796 => "10000110",
 3797 => "00000111",
 3798 => "00011100",
 3799 => "01001111",
 3800 => "11101000",
 3801 => "10000101",
 3802 => "10100010",
 3803 => "11011110",
 3804 => "01001001",
 3805 => "10101101",
 3806 => "11010011",
 3807 => "00001010",
 3808 => "01101100",
 3809 => "00100100",
 3810 => "01010000",
 3811 => "10101000",
 3812 => "00110111",
 3813 => "00110001",
 3814 => "11101111",
 3815 => "00110110",
 3816 => "10101101",
 3817 => "01111101",
 3818 => "10000011",
 3819 => "00010011",
 3820 => "00110001",
 3821 => "10000010",
 3822 => "01101100",
 3823 => "11010010",
 3824 => "10001011",
 3825 => "00001000",
 3826 => "11110110",
 3827 => "01000011",
 3828 => "00010000",
 3829 => "10111001",
 3830 => "11011000",
 3831 => "01100101",
 3832 => "00111000",
 3833 => "10101111",
 3834 => "10111100",
 3835 => "01011011",
 3836 => "00011001",
 3837 => "01001000",
 3838 => "00010001",
 3839 => "11111100",
 3840 => "10011101",
 3841 => "10111110",
 3842 => "01010010",
 3843 => "10010111",
 3844 => "11100000",
 3845 => "01100010",
 3846 => "01100001",
 3847 => "00011001",
 3848 => "01011100",
 3849 => "11000010",
 3850 => "11100011",
 3851 => "10110001",
 3852 => "11101001",
 3853 => "00000010",
 3854 => "11010011",
 3855 => "11011101",
 3856 => "10100010",
 3857 => "01000101",
 3858 => "11011000",
 3859 => "11000010",
 3860 => "01111010",
 3861 => "01000110",
 3862 => "01011100",
 3863 => "11100011",
 3864 => "10011000",
 3865 => "11000010",
 3866 => "10111011",
 3867 => "11011100",
 3868 => "01101111",
 3869 => "00010001",
 3870 => "10001000",
 3871 => "01011101",
 3872 => "11010110",
 3873 => "01010111",
 3874 => "10110010",
 3875 => "01101001",
 3876 => "10111010",
 3877 => "00101111",
 3878 => "00111111",
 3879 => "10011110",
 3880 => "10100010",
 3881 => "00110000",
 3882 => "01101011",
 3883 => "00100101",
 3884 => "10001001",
 3885 => "01000101",
 3886 => "00111110",
 3887 => "00000111",
 3888 => "00000101",
 3889 => "00011101",
 3890 => "11100010",
 3891 => "01011100",
 3892 => "10001001",
 3893 => "10110100",
 3894 => "10101100",
 3895 => "10101011",
 3896 => "11111101",
 3897 => "00110110",
 3898 => "01010000",
 3899 => "01111110",
 3900 => "01110001",
 3901 => "10100111",
 3902 => "00110110",
 3903 => "10100011",
 3904 => "01110000",
 3905 => "00011011",
 3906 => "10100001",
 3907 => "00111000",
 3908 => "11110100",
 3909 => "00110001",
 3910 => "10001110",
 3911 => "10110010",
 3912 => "00110011",
 3913 => "11010100",
 3914 => "11100010",
 3915 => "11111100",
 3916 => "01000000",
 3917 => "10000110",
 3918 => "01000010",
 3919 => "11100010",
 3920 => "11111110",
 3921 => "01000110",
 3922 => "10101101",
 3923 => "00110001",
 3924 => "10000010",
 3925 => "00000100",
 3926 => "11011000",
 3927 => "11001100",
 3928 => "11111011",
 3929 => "11100110",
 3930 => "01111110",
 3931 => "01111000",
 3932 => "11101000",
 3933 => "10100110",
 3934 => "01100000",
 3935 => "00100110",
 3936 => "00011001",
 3937 => "01110100",
 3938 => "11011000",
 3939 => "10011010",
 3940 => "00111101",
 3941 => "11110011",
 3942 => "10100000",
 3943 => "11001000",
 3944 => "10101101",
 3945 => "11010001",
 3946 => "01010001",
 3947 => "10100100",
 3948 => "11000111",
 3949 => "11110000",
 3950 => "11110000",
 3951 => "00100011",
 3952 => "01001000",
 3953 => "00001000",
 3954 => "01011000",
 3955 => "01000100",
 3956 => "10000011",
 3957 => "00001000",
 3958 => "01001010",
 3959 => "01111001",
 3960 => "10111010",
 3961 => "00110101",
 3962 => "10011001",
 3963 => "01101101",
 3964 => "10011010",
 3965 => "00010100",
 3966 => "00000001",
 3967 => "00000110",
 3968 => "10010101",
 3969 => "10101110",
 3970 => "00001000",
 3971 => "11010101",
 3972 => "11000011",
 3973 => "00100110",
 3974 => "00000011",
 3975 => "01100110",
 3976 => "11000000",
 3977 => "10111001",
 3978 => "00000011",
 3979 => "10011100",
 3980 => "01001010",
 3981 => "11001000",
 3982 => "01110000",
 3983 => "00011101",
 3984 => "10001010",
 3985 => "00000101",
 3986 => "10010001",
 3987 => "11100011",
 3988 => "10010110",
 3989 => "10011100",
 3990 => "11100000",
 3991 => "10011100",
 3992 => "11101000",
 3993 => "11101100",
 3994 => "00010111",
 3995 => "11000000",
 3996 => "11110010",
 3997 => "00110010",
 3998 => "01101011",
 3999 => "11111110",
 4000 => "10110110",
 4001 => "01101000",
 4002 => "01001001",
 4003 => "10101000",
 4004 => "10011101",
 4005 => "01111011",
 4006 => "01010000",
 4007 => "10011011",
 4008 => "01101101",
 4009 => "00011110",
 4010 => "11101100",
 4011 => "01110111",
 4012 => "10011111",
 4013 => "11000000",
 4014 => "01111011",
 4015 => "00111000",
 4016 => "11100000",
 4017 => "00011010",
 4018 => "00100011",
 4019 => "11101100",
 4020 => "10001000",
 4021 => "01010110",
 4022 => "10110110",
 4023 => "00000001",
 4024 => "11010000",
 4025 => "11100011",
 4026 => "00111011",
 4027 => "01110011",
 4028 => "10011001",
 4029 => "00001111",
 4030 => "11010000",
 4031 => "01001010",
 4032 => "01111011",
 4033 => "00111111",
 4034 => "10001111",
 4035 => "01011100",
 4036 => "10110010",
 4037 => "11100010",
 4038 => "00001111",
 4039 => "00011100",
 4040 => "00001000",
 4041 => "00101111",
 4042 => "11000001",
 4043 => "11101101",
 4044 => "01101110",
 4045 => "10011001",
 4046 => "01011001",
 4047 => "11110101",
 4048 => "00011110",
 4049 => "01101111",
 4050 => "01001101",
 4051 => "00001110",
 4052 => "00101011",
 4053 => "01101111",
 4054 => "01001100",
 4055 => "00000011",
 4056 => "00100001",
 4057 => "11101100",
 4058 => "10101001",
 4059 => "10101000",
 4060 => "01011011",
 4061 => "01010000",
 4062 => "00011111",
 4063 => "10001111",
 4064 => "01111101",
 4065 => "10110101",
 4066 => "01110000",
 4067 => "10001100",
 4068 => "01000101",
 4069 => "11011110",
 4070 => "10101000",
 4071 => "00011100",
 4072 => "00101011",
 4073 => "10100011",
 4074 => "00101101",
 4075 => "11100110",
 4076 => "00001010",
 4077 => "00100101",
 4078 => "00111001",
 4079 => "11111000",
 4080 => "11111000",
 4081 => "10111101",
 4082 => "01001001",
 4083 => "10011111",
 4084 => "01000011",
 4085 => "10010010",
 4086 => "11111001",
 4087 => "11101100",
 4088 => "11111100",
 4089 => "00100111",
 4090 => "00000011",
 4091 => "01011111",
 4092 => "01111000",
 4093 => "00010010",
 4094 => "11111000",
 4095 => "00001100",
 4096 => "01000110",
 4097 => "00000000",
 4098 => "01111011",
 4099 => "00010101",
 4100 => "10001111",
 4101 => "11011011",
 4102 => "10100011",
 4103 => "10001001",
 4104 => "01100100",
 4105 => "01000000",
 4106 => "11101001",
 4107 => "11000100",
 4108 => "01000000",
 4109 => "01110011",
 4110 => "01011010",
 4111 => "01010111",
 4112 => "00110001",
 4113 => "00011000",
 4114 => "11001110",
 4115 => "10101101",
 4116 => "01011011",
 4117 => "01011010",
 4118 => "00011100",
 4119 => "10010111",
 4120 => "10010001",
 4121 => "00010010",
 4122 => "11101000",
 4123 => "11101111",
 4124 => "00110111",
 4125 => "11111011",
 4126 => "11101000",
 4127 => "00111110",
 4128 => "10001111",
 4129 => "11010111",
 4130 => "01001010",
 4131 => "01101110",
 4132 => "01100101",
 4133 => "00010001",
 4134 => "11111111",
 4135 => "11010111",
 4136 => "01001100",
 4137 => "10001111",
 4138 => "00000101",
 4139 => "11000011",
 4140 => "01100111",
 4141 => "10110001",
 4142 => "00000101",
 4143 => "11000111",
 4144 => "01001111",
 4145 => "00010001",
 4146 => "11010010",
 4147 => "01101100",
 4148 => "10110110",
 4149 => "00100110",
 4150 => "01001000",
 4151 => "10000101",
 4152 => "10110100",
 4153 => "01100111",
 4154 => "01001101",
 4155 => "01111011",
 4156 => "00110110",
 4157 => "11010000",
 4158 => "10000101",
 4159 => "10111001",
 4160 => "10000000",
 4161 => "00101111",
 4162 => "10100100",
 4163 => "01111111",
 4164 => "10001001",
 4165 => "00111101",
 4166 => "10100000",
 4167 => "01101010",
 4168 => "00100011",
 4169 => "00010000",
 4170 => "11000000",
 4171 => "01100010",
 4172 => "01110000",
 4173 => "10110000",
 4174 => "00001001",
 4175 => "10100010",
 4176 => "01001010",
 4177 => "01011101",
 4178 => "01100101",
 4179 => "10001100",
 4180 => "01111110",
 4181 => "01010001",
 4182 => "11011110",
 4183 => "10001110",
 4184 => "10001101",
 4185 => "11011011",
 4186 => "11011100",
 4187 => "11001111",
 4188 => "01000010",
 4189 => "11010011",
 4190 => "10101101",
 4191 => "10100010",
 4192 => "00010001",
 4193 => "00110111",
 4194 => "11111100",
 4195 => "01011101",
 4196 => "01111010",
 4197 => "00100110",
 4198 => "11010100",
 4199 => "01110010",
 4200 => "10100001",
 4201 => "00100101",
 4202 => "01010100",
 4203 => "10110100",
 4204 => "10001010",
 4205 => "10101011",
 4206 => "10001011",
 4207 => "11110000",
 4208 => "00101010",
 4209 => "00000110",
 4210 => "01110000",
 4211 => "00101000",
 4212 => "01111001",
 4213 => "11011010",
 4214 => "00111101",
 4215 => "10010010",
 4216 => "10011001",
 4217 => "11101111",
 4218 => "11001100",
 4219 => "01110101",
 4220 => "01111000",
 4221 => "00101110",
 4222 => "00100000",
 4223 => "10001110",
 4224 => "11001011",
 4225 => "10101001",
 4226 => "10001001",
 4227 => "11110110",
 4228 => "01100111",
 4229 => "10011110",
 4230 => "00010010",
 4231 => "00001000",
 4232 => "11000001",
 4233 => "01001110",
 4234 => "11110101",
 4235 => "01101101",
 4236 => "01000011",
 4237 => "00100110", others => (others =>'0'));
component project_reti_logiche is 
    port (
            i_clk         : in  std_logic;
            i_start       : in  std_logic;
            i_rst         : in  std_logic;
            i_data       : in  std_logic_vector(7 downto 0); --1 byte
            o_address     : out std_logic_vector(15 downto 0); --16 bit addr: max size is 255*255 + 3 more for max x and y and thresh.
            o_done            : out std_logic;
            o_en         : out std_logic;
            o_we       : out std_logic;
            o_data            : out std_logic_vector (7 downto 0)
          );
end component project_reti_logiche;
begin 
	UUT: project_reti_logiche
	port map (
		  i_clk      	=> tb_clk,	
          i_start       => tb_start,
          i_rst      	=> tb_rst,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address, 
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
		  o_we 	=> mem_we,
          o_data    => mem_i_data
);p_CLK_GEN : process is
  begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
  end process p_CLK_GEN; 
 MEM : process(tb_clk)
   begin
    if tb_clk'event and tb_clk = '1' then
     if enable_wire = '1' then
      if mem_we = '1' then
       RAM(conv_integer(mem_address))              <= mem_i_data;
       mem_o_data                      <= mem_i_data;
      else
       mem_o_data <= RAM(conv_integer(mem_address));
      end if;
     end if;
    end if;
   end process;
test : process is
begin 
wait for 100 ns;
wait for c_CLOCK_PERIOD;
tb_rst <= '1';
wait for c_CLOCK_PERIOD;
tb_rst <= '0';
wait for c_CLOCK_PERIOD;
tb_start <= '1';
wait for c_CLOCK_PERIOD; 
tb_start <= '0';
wait until tb_done = '1';
wait until tb_done = '0';
wait until rising_edge(tb_clk);

 
assert RAM(1) = "00010000" report "FAIL high bits" severity failure;
assert RAM(0) = "10001001" report "FAIL low bits" severity failure;
assert false report "Simulation Ended!, test passed" severity failure;
end process test;
 end projecttb;