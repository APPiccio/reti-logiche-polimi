library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity project_tb is
end project_tb;
architecture projecttb of project_tb is
constant c_CLOCK_PERIOD		: time := 15 ns;
signal   tb_done		: std_logic;
signal   mem_address		: std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst		    : std_logic := '0';
signal   tb_start		: std_logic := '0';
signal   tb_clk		    : std_logic := '0';
signal   mem_o_data,mem_i_data		: std_logic_vector (7 downto 0);
signal   enable_wire  		: std_logic;
signal   mem_we		: std_logic;
type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
signal RAM: ram_type := (2 => "01100100", 3 => "01000001", 4 => "10001100",
 5 => "11100101",
 6 => "01111001",
 7 => "00110101",
 8 => "01011010",
 9 => "01001011",
 10 => "11111001",
 11 => "01101111",
 12 => "11011100",
 13 => "11001011",
 14 => "00101010",
 15 => "00101100",
 16 => "01010110",
 17 => "10001110",
 18 => "10001111",
 19 => "10101010",
 20 => "01010100",
 21 => "01101110",
 22 => "11010111",
 23 => "10000001",
 24 => "11011101",
 25 => "10001111",
 26 => "00000110",
 27 => "11101100",
 28 => "00001010",
 29 => "00110001",
 30 => "00110101",
 31 => "11110001",
 32 => "10010010",
 33 => "00110010",
 34 => "00100000",
 35 => "10010110",
 36 => "11110101",
 37 => "00010011",
 38 => "01001010",
 39 => "00101100",
 40 => "00011010",
 41 => "10000110",
 42 => "10111001",
 43 => "11000000",
 44 => "11000011",
 45 => "00000100",
 46 => "11101111",
 47 => "10011101",
 48 => "00110010",
 49 => "01010001",
 50 => "11011010",
 51 => "10110011",
 52 => "10011010",
 53 => "01101110",
 54 => "10101101",
 55 => "01101100",
 56 => "01001111",
 57 => "01110100",
 58 => "11010100",
 59 => "10110010",
 60 => "01001101",
 61 => "10011100",
 62 => "00010000",
 63 => "10101000",
 64 => "10011000",
 65 => "00011000",
 66 => "01100010",
 67 => "01101000",
 68 => "00000011",
 69 => "00000001",
 70 => "00001000",
 71 => "00001110",
 72 => "10101100",
 73 => "01000010",
 74 => "10110100",
 75 => "10110011",
 76 => "00001101",
 77 => "10011100",
 78 => "01101001",
 79 => "00010001",
 80 => "00010000",
 81 => "11010000",
 82 => "11000000",
 83 => "00001001",
 84 => "00000010",
 85 => "01000111",
 86 => "01111111",
 87 => "01001010",
 88 => "00011101",
 89 => "01101010",
 90 => "11101111",
 91 => "10001010",
 92 => "10111110",
 93 => "00011101",
 94 => "00010101",
 95 => "00000011",
 96 => "11100000",
 97 => "00011001",
 98 => "10011110",
 99 => "00110001",
 100 => "00110011",
 101 => "00010111",
 102 => "10000110",
 103 => "10011101",
 104 => "01100010",
 105 => "01010011",
 106 => "00110111",
 107 => "01001110",
 108 => "11100011",
 109 => "10110100",
 110 => "10101010",
 111 => "11110101",
 112 => "11011011",
 113 => "00010000",
 114 => "10000111",
 115 => "11111100",
 116 => "01011010",
 117 => "10001011",
 118 => "00000010",
 119 => "01100101",
 120 => "10001011",
 121 => "10010110",
 122 => "00001010",
 123 => "10111100",
 124 => "11010100",
 125 => "11011100",
 126 => "11010101",
 127 => "01010111",
 128 => "11101001",
 129 => "10011000",
 130 => "01011100",
 131 => "01001111",
 132 => "00010000",
 133 => "00110011",
 134 => "00010111",
 135 => "01011001",
 136 => "11001001",
 137 => "00101100",
 138 => "10100111",
 139 => "10110001",
 140 => "01110100",
 141 => "10111010",
 142 => "10111001",
 143 => "00001011",
 144 => "11000000",
 145 => "01101100",
 146 => "10101101",
 147 => "00111110",
 148 => "00100100",
 149 => "10010011",
 150 => "00110000",
 151 => "01001101",
 152 => "00110111",
 153 => "01010010",
 154 => "10000001",
 155 => "11000110",
 156 => "00111000",
 157 => "10100100",
 158 => "11110011",
 159 => "01111001",
 160 => "11101000",
 161 => "00010001",
 162 => "00111100",
 163 => "11000110",
 164 => "11110111",
 165 => "01011101",
 166 => "01110111",
 167 => "10000011",
 168 => "00000110",
 169 => "00001001",
 170 => "01101101",
 171 => "01000100",
 172 => "01000111",
 173 => "00010111",
 174 => "00110101",
 175 => "10111011",
 176 => "11000001",
 177 => "00001010",
 178 => "11010011",
 179 => "11011000",
 180 => "11101011",
 181 => "10010010",
 182 => "11011100",
 183 => "01111011",
 184 => "00001001",
 185 => "00001000",
 186 => "00010101",
 187 => "10011111",
 188 => "01110010",
 189 => "10110000",
 190 => "10000001",
 191 => "00000111",
 192 => "01101111",
 193 => "01100001",
 194 => "11111101",
 195 => "00100101",
 196 => "10100010",
 197 => "10111110",
 198 => "11011011",
 199 => "10010101",
 200 => "10000101",
 201 => "11110111",
 202 => "11010110",
 203 => "11001111",
 204 => "00110001",
 205 => "01011001",
 206 => "00010011",
 207 => "10111010",
 208 => "10001111",
 209 => "01000011",
 210 => "00010101",
 211 => "01111001",
 212 => "11111010",
 213 => "10101001",
 214 => "00100010",
 215 => "11010101",
 216 => "10000000",
 217 => "00100010",
 218 => "01010000",
 219 => "10000101",
 220 => "01010101",
 221 => "11001111",
 222 => "11101011",
 223 => "00010100",
 224 => "10001101",
 225 => "10110010",
 226 => "11000010",
 227 => "11001101",
 228 => "10101010",
 229 => "11000011",
 230 => "10000110",
 231 => "00100011",
 232 => "00111100",
 233 => "00010101",
 234 => "10010000",
 235 => "00001101",
 236 => "10001011",
 237 => "10000011",
 238 => "11001000",
 239 => "10101011",
 240 => "10001000",
 241 => "10101010",
 242 => "11010001",
 243 => "00001011",
 244 => "01010011",
 245 => "10110000",
 246 => "01011000",
 247 => "00101111",
 248 => "01010100",
 249 => "11000000",
 250 => "00001010",
 251 => "10010011",
 252 => "11000011",
 253 => "11000101",
 254 => "00001000",
 255 => "00000101",
 256 => "10011001",
 257 => "00110101",
 258 => "01000001",
 259 => "10001111",
 260 => "00000000",
 261 => "00101010",
 262 => "11110111",
 263 => "11001111",
 264 => "11101110",
 265 => "10110011",
 266 => "10110100",
 267 => "00011110",
 268 => "01101011",
 269 => "00111011",
 270 => "01111100",
 271 => "11010111",
 272 => "10111010",
 273 => "01011010",
 274 => "10110101",
 275 => "10000110",
 276 => "01001111",
 277 => "10101010",
 278 => "01111000",
 279 => "11110111",
 280 => "11101011",
 281 => "00001011",
 282 => "11010001",
 283 => "01001010",
 284 => "11000100",
 285 => "10011111",
 286 => "11111011",
 287 => "00101000",
 288 => "01110110",
 289 => "01101001",
 290 => "00110011",
 291 => "11001101",
 292 => "00011111",
 293 => "11001101",
 294 => "00001010",
 295 => "01111110",
 296 => "01000011",
 297 => "10001010",
 298 => "11100010",
 299 => "01101101",
 300 => "10110101",
 301 => "01000011",
 302 => "01100011",
 303 => "00011000",
 304 => "00110100",
 305 => "01101111",
 306 => "01110110",
 307 => "01110000",
 308 => "11100110",
 309 => "10111011",
 310 => "11010110",
 311 => "10010100",
 312 => "10011001",
 313 => "00101000",
 314 => "01111110",
 315 => "00001000",
 316 => "11100011",
 317 => "01010000",
 318 => "11000000",
 319 => "00100011",
 320 => "01101010",
 321 => "01001000",
 322 => "01101100",
 323 => "01001011",
 324 => "00111000",
 325 => "11000111",
 326 => "10000011",
 327 => "00100100",
 328 => "10100000",
 329 => "00010111",
 330 => "10110000",
 331 => "01000001",
 332 => "10000000",
 333 => "01100001",
 334 => "10001111",
 335 => "11110110",
 336 => "00111000",
 337 => "10000000",
 338 => "01111111",
 339 => "01100010",
 340 => "11110011",
 341 => "11100110",
 342 => "11100100",
 343 => "01011111",
 344 => "00110001",
 345 => "11000000",
 346 => "00100111",
 347 => "01110010",
 348 => "10011110",
 349 => "10000011",
 350 => "10000000",
 351 => "00010001",
 352 => "01100011",
 353 => "10111100",
 354 => "11101100",
 355 => "01000111",
 356 => "11110111",
 357 => "00001001",
 358 => "11000000",
 359 => "00100101",
 360 => "10111110",
 361 => "01100011",
 362 => "10011101",
 363 => "11101000",
 364 => "01010101",
 365 => "00100101",
 366 => "10100001",
 367 => "01000100",
 368 => "10001010",
 369 => "00101101",
 370 => "00100110",
 371 => "01101000",
 372 => "00000011",
 373 => "00011000",
 374 => "11010000",
 375 => "11010111",
 376 => "00000111",
 377 => "00000000",
 378 => "11101110",
 379 => "01011110",
 380 => "11110010",
 381 => "01011010",
 382 => "00001111",
 383 => "11101000",
 384 => "00000111",
 385 => "00001010",
 386 => "10010001",
 387 => "10010010",
 388 => "11001011",
 389 => "11011100",
 390 => "11110000",
 391 => "11111100",
 392 => "11001111",
 393 => "10010110",
 394 => "01010100",
 395 => "00010010",
 396 => "10100000",
 397 => "01000010",
 398 => "10100110",
 399 => "10110100",
 400 => "01011001",
 401 => "01001110",
 402 => "01000100",
 403 => "10001100",
 404 => "10001101",
 405 => "01100000",
 406 => "10110100",
 407 => "10000110",
 408 => "00010101",
 409 => "00100000",
 410 => "11100111",
 411 => "01110000",
 412 => "11111010",
 413 => "01010110",
 414 => "01010000",
 415 => "00110001",
 416 => "10110101",
 417 => "11011011",
 418 => "01000110",
 419 => "10010100",
 420 => "11001001",
 421 => "11100101",
 422 => "00011010",
 423 => "00000000",
 424 => "10011010",
 425 => "00111101",
 426 => "11010110",
 427 => "11111010",
 428 => "01001000",
 429 => "11000100",
 430 => "11111100",
 431 => "01110011",
 432 => "00011100",
 433 => "11111111",
 434 => "10101101",
 435 => "01111001",
 436 => "00010010",
 437 => "01000010",
 438 => "10001011",
 439 => "01100111",
 440 => "00110110",
 441 => "01100110",
 442 => "10100101",
 443 => "11100000",
 444 => "10001111",
 445 => "11110111",
 446 => "00011000",
 447 => "00011011",
 448 => "11101101",
 449 => "00110000",
 450 => "10111010",
 451 => "10111000",
 452 => "11101101",
 453 => "10100110",
 454 => "10101101",
 455 => "01101000",
 456 => "10111001",
 457 => "10110111",
 458 => "01101000",
 459 => "11101111",
 460 => "10011101",
 461 => "11110000",
 462 => "00001000",
 463 => "10001011",
 464 => "01000100",
 465 => "10011011",
 466 => "10001011",
 467 => "00011100",
 468 => "00110011",
 469 => "01000010",
 470 => "00010011",
 471 => "11100101",
 472 => "11010100",
 473 => "01010100",
 474 => "01000011",
 475 => "00101111",
 476 => "10100011",
 477 => "01111110",
 478 => "00010100",
 479 => "10111010",
 480 => "11011110",
 481 => "00001001",
 482 => "10110110",
 483 => "01100111",
 484 => "10001110",
 485 => "00101001",
 486 => "10010110",
 487 => "10110010",
 488 => "10110111",
 489 => "10000010",
 490 => "00100101",
 491 => "10000011",
 492 => "11110010",
 493 => "01010000",
 494 => "10000111",
 495 => "10110011",
 496 => "11111011",
 497 => "01111001",
 498 => "01101101",
 499 => "11100110",
 500 => "00100111",
 501 => "00101110",
 502 => "00111000",
 503 => "00110100",
 504 => "10000010",
 505 => "00001101",
 506 => "01101110",
 507 => "01001100",
 508 => "01010011",
 509 => "01001001",
 510 => "01010000",
 511 => "10011111",
 512 => "01100100",
 513 => "00010111",
 514 => "10011101",
 515 => "01011011",
 516 => "11001111",
 517 => "01001001",
 518 => "00101011",
 519 => "01111110",
 520 => "00000110",
 521 => "00010011",
 522 => "10101100",
 523 => "01000100",
 524 => "10101001",
 525 => "01101101",
 526 => "11111001",
 527 => "11001111",
 528 => "00011000",
 529 => "10011011",
 530 => "10000111",
 531 => "10100100",
 532 => "01001010",
 533 => "10001011",
 534 => "11000000",
 535 => "10001000",
 536 => "01001101",
 537 => "00101010",
 538 => "00011010",
 539 => "10010111",
 540 => "01110100",
 541 => "01111110",
 542 => "10011101",
 543 => "10011010",
 544 => "01110111",
 545 => "00011010",
 546 => "00100001",
 547 => "01110001",
 548 => "00100111",
 549 => "11010111",
 550 => "01110101",
 551 => "11110111",
 552 => "00111111",
 553 => "00001111",
 554 => "00000101",
 555 => "00011000",
 556 => "00101101",
 557 => "00101010",
 558 => "00011100",
 559 => "00110101",
 560 => "00101111",
 561 => "01010111",
 562 => "11100111",
 563 => "00001011",
 564 => "10001110",
 565 => "11010001",
 566 => "11100110",
 567 => "11010001",
 568 => "10110101",
 569 => "11001000",
 570 => "11010111",
 571 => "10011011",
 572 => "10101100",
 573 => "01001010",
 574 => "11101001",
 575 => "00011110",
 576 => "11010010",
 577 => "10000010",
 578 => "11001011",
 579 => "11111111",
 580 => "01011000",
 581 => "01001000",
 582 => "10011111",
 583 => "10111000",
 584 => "10000110",
 585 => "00100101",
 586 => "00100101",
 587 => "10110110",
 588 => "10011010",
 589 => "00100100",
 590 => "11001011",
 591 => "11000000",
 592 => "00000101",
 593 => "01110100",
 594 => "10011101",
 595 => "11100000",
 596 => "01010000",
 597 => "10011011",
 598 => "00110101",
 599 => "11101111",
 600 => "10101000",
 601 => "01001100",
 602 => "11100010",
 603 => "01110110",
 604 => "10101000",
 605 => "00110100",
 606 => "00110011",
 607 => "00000111",
 608 => "01101110",
 609 => "00010100",
 610 => "00011101",
 611 => "01010100",
 612 => "11110111",
 613 => "11000010",
 614 => "00011011",
 615 => "10001110",
 616 => "01011110",
 617 => "01100100",
 618 => "01011111",
 619 => "11000001",
 620 => "11001001",
 621 => "11101101",
 622 => "00100101",
 623 => "00001001",
 624 => "01110101",
 625 => "01111110",
 626 => "11100000",
 627 => "11100110",
 628 => "10101011",
 629 => "00001100",
 630 => "00010100",
 631 => "01101111",
 632 => "01010011",
 633 => "11101110",
 634 => "00000001",
 635 => "10110111",
 636 => "01111000",
 637 => "10111100",
 638 => "01100110",
 639 => "01101001",
 640 => "00100011",
 641 => "01111110",
 642 => "00111100",
 643 => "01101101",
 644 => "00101000",
 645 => "10001110",
 646 => "00100110",
 647 => "11100000",
 648 => "11000001",
 649 => "11101001",
 650 => "00101100",
 651 => "10011010",
 652 => "00111101",
 653 => "10111000",
 654 => "10000011",
 655 => "11010100",
 656 => "00001010",
 657 => "00010010",
 658 => "11100110",
 659 => "01010110",
 660 => "00000101",
 661 => "10000010",
 662 => "01100000",
 663 => "01100110",
 664 => "10100101",
 665 => "01011011",
 666 => "11110011",
 667 => "11101100",
 668 => "10001011",
 669 => "11010101",
 670 => "00000001",
 671 => "10011000",
 672 => "10010001",
 673 => "01001000",
 674 => "11100101",
 675 => "01111010",
 676 => "01000111",
 677 => "01110111",
 678 => "01110001",
 679 => "10101001",
 680 => "10100010",
 681 => "01100011",
 682 => "10100101",
 683 => "01111010",
 684 => "00111111",
 685 => "11001101",
 686 => "01000001",
 687 => "11011101",
 688 => "00000111",
 689 => "11111000",
 690 => "10100011",
 691 => "00111100",
 692 => "10100001",
 693 => "01010000",
 694 => "01010110",
 695 => "10100101",
 696 => "10101010",
 697 => "00111011",
 698 => "10000111",
 699 => "00101110",
 700 => "00000110",
 701 => "10100100",
 702 => "01001100",
 703 => "10011110",
 704 => "00111010",
 705 => "01110011",
 706 => "00111001",
 707 => "01001100",
 708 => "00101000",
 709 => "00011110",
 710 => "11110111",
 711 => "11110001",
 712 => "11110010",
 713 => "00100111",
 714 => "11111111",
 715 => "10001110",
 716 => "00110000",
 717 => "00011110",
 718 => "00000000",
 719 => "11110001",
 720 => "11111001",
 721 => "01101011",
 722 => "11010000",
 723 => "11110100",
 724 => "11101000",
 725 => "11111000",
 726 => "10001001",
 727 => "01110000",
 728 => "11001100",
 729 => "00100011",
 730 => "11100001",
 731 => "00010001",
 732 => "10111100",
 733 => "01111111",
 734 => "10000010",
 735 => "00101110",
 736 => "10111101",
 737 => "01111010",
 738 => "00110110",
 739 => "01110101",
 740 => "10010001",
 741 => "01001101",
 742 => "01101010",
 743 => "10110100",
 744 => "00000100",
 745 => "10110101",
 746 => "10001101",
 747 => "10011101",
 748 => "01001101",
 749 => "10100000",
 750 => "11110011",
 751 => "01000000",
 752 => "10000011",
 753 => "10110100",
 754 => "01011111",
 755 => "10011100",
 756 => "11000000",
 757 => "10110100",
 758 => "11110011",
 759 => "11010011",
 760 => "01110110",
 761 => "00100011",
 762 => "11111011",
 763 => "00011101",
 764 => "11001111",
 765 => "10011001",
 766 => "11000010",
 767 => "10101010",
 768 => "11001000",
 769 => "10110111",
 770 => "10100110",
 771 => "11101000",
 772 => "10100101",
 773 => "00000100",
 774 => "11100110",
 775 => "01011111",
 776 => "10110010",
 777 => "11010101",
 778 => "00110011",
 779 => "10011111",
 780 => "11011111",
 781 => "11111101",
 782 => "01111110",
 783 => "10101011",
 784 => "00101101",
 785 => "00010011",
 786 => "01100000",
 787 => "00000001",
 788 => "10101000",
 789 => "01011010",
 790 => "10111110",
 791 => "01000110",
 792 => "01101010",
 793 => "01110111",
 794 => "00111001",
 795 => "01000011",
 796 => "10111111",
 797 => "00111101",
 798 => "01111001",
 799 => "10101001",
 800 => "10011111",
 801 => "00110011",
 802 => "00110111",
 803 => "00011101",
 804 => "00111111",
 805 => "00100000",
 806 => "00000111",
 807 => "11111010",
 808 => "10011010",
 809 => "00101111",
 810 => "01111001",
 811 => "11001001",
 812 => "11001100",
 813 => "10101111",
 814 => "10100011",
 815 => "00101000",
 816 => "01001000",
 817 => "01111001",
 818 => "01110101",
 819 => "11101010",
 820 => "00100111",
 821 => "00110011",
 822 => "10101000",
 823 => "10010101",
 824 => "01010111",
 825 => "11000100",
 826 => "11101100",
 827 => "11111100",
 828 => "11100111",
 829 => "10001111",
 830 => "00001110",
 831 => "00110101",
 832 => "01111101",
 833 => "01011010",
 834 => "01110001",
 835 => "00100000",
 836 => "11110011",
 837 => "10001001",
 838 => "10100111",
 839 => "11100010",
 840 => "11111110",
 841 => "11100101",
 842 => "00101111",
 843 => "00111110",
 844 => "11011001",
 845 => "00010010",
 846 => "00111010",
 847 => "10100100",
 848 => "01010101",
 849 => "11010101",
 850 => "11100010",
 851 => "10110010",
 852 => "01100100",
 853 => "01111011",
 854 => "00010101",
 855 => "10110010",
 856 => "01001011",
 857 => "11100110",
 858 => "00000011",
 859 => "10100010",
 860 => "00111101",
 861 => "01111010",
 862 => "00001011",
 863 => "10000000",
 864 => "00000001",
 865 => "00101010",
 866 => "10110000",
 867 => "01111101",
 868 => "00010011",
 869 => "00101010",
 870 => "00011010",
 871 => "00110011",
 872 => "00110101",
 873 => "11111000",
 874 => "00101110",
 875 => "00000101",
 876 => "10001010",
 877 => "00000011",
 878 => "00001101",
 879 => "11110000",
 880 => "10010110",
 881 => "10110000",
 882 => "10000111",
 883 => "01100000",
 884 => "11100011",
 885 => "00100010",
 886 => "11100010",
 887 => "10111101",
 888 => "00010101",
 889 => "00110001",
 890 => "10001101",
 891 => "11001011",
 892 => "10111100",
 893 => "10101001",
 894 => "00111111",
 895 => "10110011",
 896 => "10010000",
 897 => "00111010",
 898 => "01001111",
 899 => "11010100",
 900 => "00111000",
 901 => "11001000",
 902 => "11110001",
 903 => "11010100",
 904 => "10101101",
 905 => "11000010",
 906 => "11000101",
 907 => "11100110",
 908 => "00111110",
 909 => "01001110",
 910 => "00110100",
 911 => "01001100",
 912 => "01011101",
 913 => "11011110",
 914 => "00111110",
 915 => "10100011",
 916 => "00101110",
 917 => "01000100",
 918 => "11111011",
 919 => "01101000",
 920 => "11110010",
 921 => "00111111",
 922 => "01011100",
 923 => "11101101",
 924 => "00110100",
 925 => "10000111",
 926 => "00111000",
 927 => "10100001",
 928 => "11001010",
 929 => "10101011",
 930 => "10001000",
 931 => "00100110",
 932 => "10011000",
 933 => "01101000",
 934 => "10001100",
 935 => "10001000",
 936 => "10001111",
 937 => "01111010",
 938 => "11100010",
 939 => "11000011",
 940 => "11000001",
 941 => "11111101",
 942 => "00001111",
 943 => "00100000",
 944 => "10010010",
 945 => "10011001",
 946 => "01110001",
 947 => "01010000",
 948 => "10000100",
 949 => "10010000",
 950 => "11111001",
 951 => "00110111",
 952 => "00000101",
 953 => "10110010",
 954 => "11001101",
 955 => "01110110",
 956 => "01100001",
 957 => "01111101",
 958 => "10010101",
 959 => "10111111",
 960 => "01010101",
 961 => "11110001",
 962 => "10001111",
 963 => "11111110",
 964 => "10100001",
 965 => "00000011",
 966 => "00100011",
 967 => "10010110",
 968 => "10111100",
 969 => "00011101",
 970 => "11110111",
 971 => "01110001",
 972 => "11000110",
 973 => "10101010",
 974 => "01010111",
 975 => "10101000",
 976 => "00101000",
 977 => "11001001",
 978 => "00100001",
 979 => "10000001",
 980 => "10011100",
 981 => "10000110",
 982 => "10100101",
 983 => "01110001",
 984 => "11000111",
 985 => "00000111",
 986 => "01010010",
 987 => "00010110",
 988 => "11010100",
 989 => "01011110",
 990 => "00111010",
 991 => "01101000",
 992 => "00000100",
 993 => "11110011",
 994 => "11001100",
 995 => "11111010",
 996 => "10101011",
 997 => "00000101",
 998 => "00001011",
 999 => "01110010",
 1000 => "10110111",
 1001 => "10101110",
 1002 => "01010111",
 1003 => "11101111",
 1004 => "01100110",
 1005 => "10001010",
 1006 => "11100110",
 1007 => "01010001",
 1008 => "10100101",
 1009 => "10001000",
 1010 => "10111110",
 1011 => "10010100",
 1012 => "10000011",
 1013 => "01011111",
 1014 => "10110010",
 1015 => "10111110",
 1016 => "00101111",
 1017 => "10100010",
 1018 => "01110100",
 1019 => "11100011",
 1020 => "00010001",
 1021 => "01000100",
 1022 => "00101010",
 1023 => "10011010",
 1024 => "10001101",
 1025 => "01100101",
 1026 => "10111111",
 1027 => "10011001",
 1028 => "11001011",
 1029 => "10100111",
 1030 => "10001011",
 1031 => "00100101",
 1032 => "00100011",
 1033 => "10011010",
 1034 => "00011101",
 1035 => "00111010",
 1036 => "00010001",
 1037 => "11101100",
 1038 => "01011011",
 1039 => "11100101",
 1040 => "10111011",
 1041 => "00001111",
 1042 => "10100000",
 1043 => "00011010",
 1044 => "11011100",
 1045 => "10011010",
 1046 => "01111010",
 1047 => "00100110",
 1048 => "01100100",
 1049 => "11101010",
 1050 => "01110001",
 1051 => "11100101",
 1052 => "01110000",
 1053 => "00110100",
 1054 => "11100010",
 1055 => "10001110",
 1056 => "01101000",
 1057 => "11000111",
 1058 => "01101000",
 1059 => "11000111",
 1060 => "00100100",
 1061 => "10110001",
 1062 => "00101100",
 1063 => "11101100",
 1064 => "00101010",
 1065 => "00100001",
 1066 => "01111100",
 1067 => "00011010",
 1068 => "11010010",
 1069 => "00111010",
 1070 => "11100011",
 1071 => "10001100",
 1072 => "10001000",
 1073 => "11101011",
 1074 => "01110001",
 1075 => "10001110",
 1076 => "00010110",
 1077 => "11110111",
 1078 => "00101001",
 1079 => "10010001",
 1080 => "11010000",
 1081 => "10111001",
 1082 => "11110111",
 1083 => "00101101",
 1084 => "00100110",
 1085 => "00011010",
 1086 => "10011010",
 1087 => "00110101",
 1088 => "00010010",
 1089 => "10100100",
 1090 => "01001010",
 1091 => "01010001",
 1092 => "01101100",
 1093 => "10011010",
 1094 => "00101111",
 1095 => "01101110",
 1096 => "11111111",
 1097 => "10111111",
 1098 => "00001100",
 1099 => "01011011",
 1100 => "10100000",
 1101 => "00001110",
 1102 => "10100100",
 1103 => "00010011",
 1104 => "10110110",
 1105 => "11010011",
 1106 => "01101111",
 1107 => "00001110",
 1108 => "00011110",
 1109 => "01101100",
 1110 => "10001110",
 1111 => "11000001",
 1112 => "01011100",
 1113 => "01000111",
 1114 => "00000000",
 1115 => "00011101",
 1116 => "01111101",
 1117 => "01100110",
 1118 => "01100011",
 1119 => "01111111",
 1120 => "11111100",
 1121 => "11110111",
 1122 => "10100110",
 1123 => "00000101",
 1124 => "11100100",
 1125 => "10110011",
 1126 => "00100011",
 1127 => "01000000",
 1128 => "10100110",
 1129 => "10101000",
 1130 => "01101101",
 1131 => "00110100",
 1132 => "00011010",
 1133 => "11010111",
 1134 => "01010110",
 1135 => "01100000",
 1136 => "00010111",
 1137 => "00001111",
 1138 => "00101100",
 1139 => "00001101",
 1140 => "01101011",
 1141 => "00001011",
 1142 => "10111001",
 1143 => "01110111",
 1144 => "00010000",
 1145 => "11000001",
 1146 => "10011110",
 1147 => "11111010",
 1148 => "10000101",
 1149 => "00100110",
 1150 => "01001000",
 1151 => "01010011",
 1152 => "00111101",
 1153 => "10011010",
 1154 => "11000110",
 1155 => "10100111",
 1156 => "10111111",
 1157 => "11001011",
 1158 => "00110010",
 1159 => "10101101",
 1160 => "01010001",
 1161 => "00010000",
 1162 => "01111111",
 1163 => "00101101",
 1164 => "11110100",
 1165 => "11001100",
 1166 => "10000111",
 1167 => "10000000",
 1168 => "10001111",
 1169 => "00010011",
 1170 => "00110010",
 1171 => "01101010",
 1172 => "11000000",
 1173 => "10011111",
 1174 => "11000000",
 1175 => "00110101",
 1176 => "10110001",
 1177 => "01000100",
 1178 => "11111010",
 1179 => "01110011",
 1180 => "00001010",
 1181 => "11011101",
 1182 => "00011101",
 1183 => "00000100",
 1184 => "11011011",
 1185 => "11011111",
 1186 => "11010011",
 1187 => "10100000",
 1188 => "10010110",
 1189 => "00111001",
 1190 => "00011000",
 1191 => "00001010",
 1192 => "11000111",
 1193 => "00000100",
 1194 => "11010001",
 1195 => "01110101",
 1196 => "01101010",
 1197 => "11001010",
 1198 => "11011111",
 1199 => "00001000",
 1200 => "01100010",
 1201 => "00101000",
 1202 => "11010110",
 1203 => "01001011",
 1204 => "00110111",
 1205 => "01010110",
 1206 => "10000011",
 1207 => "01011011",
 1208 => "01010001",
 1209 => "01000101",
 1210 => "11111111",
 1211 => "00010011",
 1212 => "01100010",
 1213 => "01111000",
 1214 => "01101111",
 1215 => "01110101",
 1216 => "00100011",
 1217 => "00100001",
 1218 => "11110100",
 1219 => "10111010",
 1220 => "01100110",
 1221 => "10100110",
 1222 => "01000000",
 1223 => "00010101",
 1224 => "11010110",
 1225 => "11000110",
 1226 => "11010011",
 1227 => "01010111",
 1228 => "00111110",
 1229 => "11100001",
 1230 => "01100001",
 1231 => "11010010",
 1232 => "00110100",
 1233 => "01011000",
 1234 => "11100110",
 1235 => "10000011",
 1236 => "10001101",
 1237 => "10110111",
 1238 => "00101000",
 1239 => "10101010",
 1240 => "10110001",
 1241 => "00101010",
 1242 => "00100101",
 1243 => "00111100",
 1244 => "00111011",
 1245 => "01000100",
 1246 => "01001100",
 1247 => "01110110",
 1248 => "00110011",
 1249 => "00110000",
 1250 => "00101000",
 1251 => "10000011",
 1252 => "11101011",
 1253 => "00001000",
 1254 => "00101011",
 1255 => "11010000",
 1256 => "11111011",
 1257 => "11000101",
 1258 => "11000011",
 1259 => "00011001",
 1260 => "00110101",
 1261 => "11100100",
 1262 => "00010100",
 1263 => "10111100",
 1264 => "00010010",
 1265 => "01101110",
 1266 => "00101100",
 1267 => "11010100",
 1268 => "01010110",
 1269 => "00110101",
 1270 => "10111010",
 1271 => "10111001",
 1272 => "10101111",
 1273 => "00011110",
 1274 => "00001011",
 1275 => "10111111",
 1276 => "00100000",
 1277 => "11110101",
 1278 => "11000110",
 1279 => "10000000",
 1280 => "00011110",
 1281 => "00110110",
 1282 => "11001110",
 1283 => "11101110",
 1284 => "00101001",
 1285 => "11100100",
 1286 => "01001111",
 1287 => "00010011",
 1288 => "10011001",
 1289 => "10111001",
 1290 => "11001101",
 1291 => "10110110",
 1292 => "01011010",
 1293 => "00110110",
 1294 => "00000110",
 1295 => "11001110",
 1296 => "01111001",
 1297 => "01000100",
 1298 => "00110110",
 1299 => "10110110",
 1300 => "11010001",
 1301 => "01000000",
 1302 => "10010101",
 1303 => "00110101",
 1304 => "01000001",
 1305 => "11111111",
 1306 => "00011111",
 1307 => "11000100",
 1308 => "01100110",
 1309 => "10001100",
 1310 => "10100111",
 1311 => "10110000",
 1312 => "01010110",
 1313 => "11101110",
 1314 => "10100011",
 1315 => "00101011",
 1316 => "00110011",
 1317 => "01101010",
 1318 => "01110101",
 1319 => "01010000",
 1320 => "11010010",
 1321 => "11000101",
 1322 => "10011010",
 1323 => "00010111",
 1324 => "00111101",
 1325 => "00000111",
 1326 => "00001111",
 1327 => "00011111",
 1328 => "11000110",
 1329 => "11011110",
 1330 => "11010111",
 1331 => "01110011",
 1332 => "11110100",
 1333 => "01010110",
 1334 => "01100111",
 1335 => "00001001",
 1336 => "01001110",
 1337 => "11011110",
 1338 => "00111001",
 1339 => "00101111",
 1340 => "11010101",
 1341 => "10101010",
 1342 => "11011011",
 1343 => "11001010",
 1344 => "00110000",
 1345 => "00111000",
 1346 => "10000001",
 1347 => "10100100",
 1348 => "10001011",
 1349 => "01110110",
 1350 => "00001100",
 1351 => "00000001",
 1352 => "01001100",
 1353 => "01101111",
 1354 => "10000100",
 1355 => "11100100",
 1356 => "01111000",
 1357 => "10010001",
 1358 => "10011001",
 1359 => "00101010",
 1360 => "10000000",
 1361 => "01111001",
 1362 => "10010100",
 1363 => "00001011",
 1364 => "11101000",
 1365 => "10010000",
 1366 => "10010000",
 1367 => "01111000",
 1368 => "10110101",
 1369 => "00101001",
 1370 => "01101111",
 1371 => "10100101",
 1372 => "00111111",
 1373 => "00011011",
 1374 => "11100000",
 1375 => "11010110",
 1376 => "11001111",
 1377 => "01001001",
 1378 => "10101011",
 1379 => "11101001",
 1380 => "00011010",
 1381 => "11000011",
 1382 => "11011010",
 1383 => "01010010",
 1384 => "10100000",
 1385 => "11001101",
 1386 => "11100100",
 1387 => "10011101",
 1388 => "10011111",
 1389 => "00001110",
 1390 => "01000101",
 1391 => "01011101",
 1392 => "01001110",
 1393 => "01010100",
 1394 => "00001101",
 1395 => "00111001",
 1396 => "10110010",
 1397 => "10101011",
 1398 => "00010110",
 1399 => "11100011",
 1400 => "01111010",
 1401 => "11100100",
 1402 => "10001011",
 1403 => "00110100",
 1404 => "01000001",
 1405 => "10111100",
 1406 => "00100001",
 1407 => "10000000",
 1408 => "01011111",
 1409 => "01011001",
 1410 => "00010011",
 1411 => "00110111",
 1412 => "01011110",
 1413 => "10110010",
 1414 => "00101101",
 1415 => "11101110",
 1416 => "11111100",
 1417 => "11001000",
 1418 => "11111010",
 1419 => "11000010",
 1420 => "11011010",
 1421 => "01100001",
 1422 => "10001101",
 1423 => "01010110",
 1424 => "11110010",
 1425 => "11100010",
 1426 => "01100111",
 1427 => "10010100",
 1428 => "11001101",
 1429 => "11010000",
 1430 => "00110110",
 1431 => "00100101",
 1432 => "11011101",
 1433 => "11010101",
 1434 => "01111001",
 1435 => "10100100",
 1436 => "10010001",
 1437 => "01001001",
 1438 => "01000010",
 1439 => "00001000",
 1440 => "10010110",
 1441 => "00011010",
 1442 => "00111010",
 1443 => "10110111",
 1444 => "11101101",
 1445 => "10000011",
 1446 => "11100101",
 1447 => "01000010",
 1448 => "01000100",
 1449 => "10101001",
 1450 => "11101011",
 1451 => "00111111",
 1452 => "10100000",
 1453 => "11101010",
 1454 => "00001110",
 1455 => "00101010",
 1456 => "01111010",
 1457 => "11011101",
 1458 => "01000111",
 1459 => "00111011",
 1460 => "10001001",
 1461 => "10000110",
 1462 => "00010101",
 1463 => "10110011",
 1464 => "00001110",
 1465 => "00100011",
 1466 => "01001001",
 1467 => "10011111",
 1468 => "10111001",
 1469 => "01101111",
 1470 => "00011100",
 1471 => "01110111",
 1472 => "00101010",
 1473 => "11000010",
 1474 => "11101100",
 1475 => "10000001",
 1476 => "01100011",
 1477 => "10001010",
 1478 => "00110001",
 1479 => "00000110",
 1480 => "00011101",
 1481 => "01010100",
 1482 => "11101110",
 1483 => "00100110",
 1484 => "10001001",
 1485 => "01100100",
 1486 => "11010111",
 1487 => "11111000",
 1488 => "00000111",
 1489 => "11011100",
 1490 => "00010111",
 1491 => "01101101",
 1492 => "11111001",
 1493 => "00111001",
 1494 => "01011110",
 1495 => "01101111",
 1496 => "00101110",
 1497 => "00000000",
 1498 => "10011011",
 1499 => "01010110",
 1500 => "01010101",
 1501 => "11111001",
 1502 => "00111001",
 1503 => "10010011",
 1504 => "01000101",
 1505 => "01011111",
 1506 => "11110110",
 1507 => "10110010",
 1508 => "11101100",
 1509 => "01010010",
 1510 => "00101000",
 1511 => "01010100",
 1512 => "10111011",
 1513 => "11001101",
 1514 => "01000011",
 1515 => "01011010",
 1516 => "11100110",
 1517 => "10101101",
 1518 => "01011010",
 1519 => "10010001",
 1520 => "00001101",
 1521 => "10101111",
 1522 => "00100001",
 1523 => "00110110",
 1524 => "10011001",
 1525 => "00101111",
 1526 => "10001110",
 1527 => "01111011",
 1528 => "00100100",
 1529 => "00010001",
 1530 => "11111101",
 1531 => "00100111",
 1532 => "10101001",
 1533 => "10111001",
 1534 => "00110010",
 1535 => "10110010",
 1536 => "01101111",
 1537 => "00101100",
 1538 => "01101100",
 1539 => "01011110",
 1540 => "01110100",
 1541 => "10001011",
 1542 => "10010111",
 1543 => "01000111",
 1544 => "01001110",
 1545 => "11001111",
 1546 => "00100010",
 1547 => "01011111",
 1548 => "01011100",
 1549 => "00101010",
 1550 => "11001100",
 1551 => "01010011",
 1552 => "00111011",
 1553 => "01000000",
 1554 => "01000001",
 1555 => "00001110",
 1556 => "01110101",
 1557 => "10110100",
 1558 => "10000000",
 1559 => "01011110",
 1560 => "10001001",
 1561 => "00101000",
 1562 => "11001000",
 1563 => "01100001",
 1564 => "00011001",
 1565 => "11001001",
 1566 => "10000101",
 1567 => "10111000",
 1568 => "00100111",
 1569 => "00110000",
 1570 => "01000000",
 1571 => "00011001",
 1572 => "11011011",
 1573 => "00111111",
 1574 => "10010011",
 1575 => "11010100",
 1576 => "10011111",
 1577 => "00001100",
 1578 => "01111010",
 1579 => "01110001",
 1580 => "01001100",
 1581 => "10101100",
 1582 => "01101101",
 1583 => "01111001",
 1584 => "00111000",
 1585 => "01110010",
 1586 => "00110000",
 1587 => "10011110",
 1588 => "01000000",
 1589 => "10011100",
 1590 => "00011010",
 1591 => "10001100",
 1592 => "10011010",
 1593 => "01100001",
 1594 => "10011011",
 1595 => "00010101",
 1596 => "00110011",
 1597 => "00101111",
 1598 => "11110001",
 1599 => "11010101",
 1600 => "10111100",
 1601 => "10010000",
 1602 => "00011011",
 1603 => "11001001",
 1604 => "11010010",
 1605 => "10101010",
 1606 => "10001101",
 1607 => "11010101",
 1608 => "10000011",
 1609 => "11111100",
 1610 => "11100100",
 1611 => "01010010",
 1612 => "10000111",
 1613 => "11001011",
 1614 => "01001010",
 1615 => "01000101",
 1616 => "00000101",
 1617 => "01001101",
 1618 => "01101010",
 1619 => "00110001",
 1620 => "00100110",
 1621 => "01101110",
 1622 => "11101111",
 1623 => "00000110",
 1624 => "01100000",
 1625 => "10101101",
 1626 => "11001010",
 1627 => "11011010",
 1628 => "10110101",
 1629 => "01111011",
 1630 => "10001001",
 1631 => "01111000",
 1632 => "11111101",
 1633 => "10110011",
 1634 => "01000011",
 1635 => "01001001",
 1636 => "11100111",
 1637 => "11010010",
 1638 => "01010110",
 1639 => "11110111",
 1640 => "11110111",
 1641 => "11110101",
 1642 => "01110001",
 1643 => "11010110",
 1644 => "11101001",
 1645 => "11001101",
 1646 => "11110100",
 1647 => "11100100",
 1648 => "11101001",
 1649 => "01011011",
 1650 => "01001111",
 1651 => "10010001",
 1652 => "10111100",
 1653 => "01100101",
 1654 => "11100101",
 1655 => "11001001",
 1656 => "11001110",
 1657 => "01111010",
 1658 => "10101110",
 1659 => "10000011",
 1660 => "10010010",
 1661 => "10111001",
 1662 => "11001111",
 1663 => "00000101",
 1664 => "01111001",
 1665 => "10000100",
 1666 => "00001000",
 1667 => "11101110",
 1668 => "10010001",
 1669 => "01111100",
 1670 => "11101010",
 1671 => "11010100",
 1672 => "01100010",
 1673 => "01011110",
 1674 => "00010101",
 1675 => "01011011",
 1676 => "00001000",
 1677 => "11111011",
 1678 => "11001001",
 1679 => "10011110",
 1680 => "00001011",
 1681 => "10101000",
 1682 => "11111011",
 1683 => "00011100",
 1684 => "10110110",
 1685 => "10101011",
 1686 => "10010011",
 1687 => "00111011",
 1688 => "10011111",
 1689 => "10000111",
 1690 => "11110000",
 1691 => "11001101",
 1692 => "01010000",
 1693 => "00000101",
 1694 => "01000001",
 1695 => "11000101",
 1696 => "00001110",
 1697 => "01101100",
 1698 => "10100110",
 1699 => "10001100",
 1700 => "11000100",
 1701 => "10110101",
 1702 => "11000001",
 1703 => "10101001",
 1704 => "00101001",
 1705 => "01110011",
 1706 => "10001110",
 1707 => "11110101",
 1708 => "11011110",
 1709 => "10111011",
 1710 => "10001101",
 1711 => "00100110",
 1712 => "10110011",
 1713 => "01010110",
 1714 => "00011101",
 1715 => "00001011",
 1716 => "00111000",
 1717 => "11011000",
 1718 => "01100001",
 1719 => "00001110",
 1720 => "00111010",
 1721 => "01101010",
 1722 => "10110100",
 1723 => "11010100",
 1724 => "10111100",
 1725 => "01111010",
 1726 => "01110101",
 1727 => "00100000",
 1728 => "01110001",
 1729 => "10010100",
 1730 => "00101111",
 1731 => "10100100",
 1732 => "00111111",
 1733 => "11100000",
 1734 => "11010001",
 1735 => "11011000",
 1736 => "00101100",
 1737 => "00001010",
 1738 => "01010110",
 1739 => "01111000",
 1740 => "10101100",
 1741 => "10100010",
 1742 => "11010100",
 1743 => "01001001",
 1744 => "10100000",
 1745 => "00101001",
 1746 => "00101011",
 1747 => "00001010",
 1748 => "01010110",
 1749 => "10111101",
 1750 => "01111111",
 1751 => "10000100",
 1752 => "11010101",
 1753 => "10110111",
 1754 => "00001011",
 1755 => "00011111",
 1756 => "10101010",
 1757 => "11011011",
 1758 => "11011001",
 1759 => "00000101",
 1760 => "11101110",
 1761 => "01110100",
 1762 => "01000100",
 1763 => "11010111",
 1764 => "10001001",
 1765 => "00100011",
 1766 => "01111100",
 1767 => "11100111",
 1768 => "01100111",
 1769 => "11001001",
 1770 => "10111011",
 1771 => "01100000",
 1772 => "10110101",
 1773 => "01110001",
 1774 => "10100010",
 1775 => "00111010",
 1776 => "11110000",
 1777 => "10111110",
 1778 => "00111110",
 1779 => "11101110",
 1780 => "11011010",
 1781 => "01100011",
 1782 => "11000001",
 1783 => "01000110",
 1784 => "00101000",
 1785 => "10111000",
 1786 => "00001011",
 1787 => "11110011",
 1788 => "01001101",
 1789 => "11101110",
 1790 => "00001010",
 1791 => "11101101",
 1792 => "10110001",
 1793 => "10000111",
 1794 => "00100000",
 1795 => "10010100",
 1796 => "11110001",
 1797 => "11100101",
 1798 => "00000101",
 1799 => "01101101",
 1800 => "11100110",
 1801 => "01010100",
 1802 => "01000010",
 1803 => "01010001",
 1804 => "11100111",
 1805 => "11011100",
 1806 => "10000001",
 1807 => "10110101",
 1808 => "11101110",
 1809 => "11110100",
 1810 => "00111001",
 1811 => "10101000",
 1812 => "10010110",
 1813 => "10001011",
 1814 => "10000011",
 1815 => "11010011",
 1816 => "00010010",
 1817 => "01011110",
 1818 => "00100011",
 1819 => "01000010",
 1820 => "11110000",
 1821 => "11100011",
 1822 => "11111010",
 1823 => "00011101",
 1824 => "01111101",
 1825 => "11010110",
 1826 => "01111110",
 1827 => "11010011",
 1828 => "11101111",
 1829 => "01100011",
 1830 => "00111000",
 1831 => "10010010",
 1832 => "11110000",
 1833 => "01111011",
 1834 => "11100001",
 1835 => "10000111",
 1836 => "11000100",
 1837 => "11001101",
 1838 => "11110111",
 1839 => "10011011",
 1840 => "10010011",
 1841 => "10101101",
 1842 => "11011000",
 1843 => "00001000",
 1844 => "10000111",
 1845 => "10111111",
 1846 => "01011000",
 1847 => "10001011",
 1848 => "00010011",
 1849 => "00000010",
 1850 => "01111110",
 1851 => "11001111",
 1852 => "00111010",
 1853 => "10011000",
 1854 => "00011111",
 1855 => "10111111",
 1856 => "00001010",
 1857 => "01101011",
 1858 => "11110111",
 1859 => "10101100",
 1860 => "00000010",
 1861 => "00110001",
 1862 => "10001110",
 1863 => "10110101",
 1864 => "01011001",
 1865 => "11111001",
 1866 => "10000100",
 1867 => "11101001",
 1868 => "00010010",
 1869 => "10101111",
 1870 => "10111101",
 1871 => "00001010",
 1872 => "00011001",
 1873 => "00000111",
 1874 => "01011111",
 1875 => "00000110",
 1876 => "01100010",
 1877 => "00001100",
 1878 => "00011110",
 1879 => "11110010",
 1880 => "10101001",
 1881 => "00100000",
 1882 => "00010010",
 1883 => "10011001",
 1884 => "01111111",
 1885 => "00001110",
 1886 => "01001100",
 1887 => "00011110",
 1888 => "00101011",
 1889 => "11001001",
 1890 => "00011100",
 1891 => "11100010",
 1892 => "10010100",
 1893 => "01011010",
 1894 => "11110111",
 1895 => "11111011",
 1896 => "10110010",
 1897 => "10111011",
 1898 => "10110100",
 1899 => "00101100",
 1900 => "10000101",
 1901 => "00111100",
 1902 => "00011111",
 1903 => "11111100",
 1904 => "10000100",
 1905 => "10111100",
 1906 => "10010101",
 1907 => "10000110",
 1908 => "10011100",
 1909 => "01101000",
 1910 => "00010001",
 1911 => "10011000",
 1912 => "01000110",
 1913 => "01011110",
 1914 => "10000010",
 1915 => "11011010",
 1916 => "11110110",
 1917 => "11111010",
 1918 => "10000001",
 1919 => "11001011",
 1920 => "00000111",
 1921 => "10001101",
 1922 => "00010110",
 1923 => "00110111",
 1924 => "11011010",
 1925 => "00011011",
 1926 => "00111000",
 1927 => "01001101",
 1928 => "01110100",
 1929 => "11001110",
 1930 => "11110100",
 1931 => "00001000",
 1932 => "10011101",
 1933 => "10000000",
 1934 => "10010001",
 1935 => "01010101",
 1936 => "00001111",
 1937 => "10000011",
 1938 => "00011101",
 1939 => "01011101",
 1940 => "00000101",
 1941 => "11101000",
 1942 => "00000111",
 1943 => "10010011",
 1944 => "10100110",
 1945 => "00001011",
 1946 => "01111101",
 1947 => "01001000",
 1948 => "10010101",
 1949 => "10000100",
 1950 => "11110111",
 1951 => "10110011",
 1952 => "00011010",
 1953 => "10001001",
 1954 => "10100100",
 1955 => "11000011",
 1956 => "00010101",
 1957 => "11110010",
 1958 => "01010111",
 1959 => "00001001",
 1960 => "11010101",
 1961 => "00000000",
 1962 => "10111011",
 1963 => "11011110",
 1964 => "00000011",
 1965 => "10011010",
 1966 => "11001011",
 1967 => "10100000",
 1968 => "01101001",
 1969 => "01100010",
 1970 => "10101010",
 1971 => "00111111",
 1972 => "10111110",
 1973 => "01001110",
 1974 => "00000101",
 1975 => "10110011",
 1976 => "10011101",
 1977 => "10001111",
 1978 => "10000010",
 1979 => "01100101",
 1980 => "01101000",
 1981 => "10101011",
 1982 => "01001110",
 1983 => "10111000",
 1984 => "10101000",
 1985 => "10110010",
 1986 => "01100001",
 1987 => "01111111",
 1988 => "00010010",
 1989 => "11011111",
 1990 => "10111000",
 1991 => "00111101",
 1992 => "01000101",
 1993 => "00000101",
 1994 => "00000001",
 1995 => "10000111",
 1996 => "11000101",
 1997 => "00110101",
 1998 => "11101001",
 1999 => "01000101",
 2000 => "00110000",
 2001 => "10100101",
 2002 => "11000011",
 2003 => "10010110",
 2004 => "11111001",
 2005 => "10110100",
 2006 => "01101010",
 2007 => "01110000",
 2008 => "10111001",
 2009 => "01010101",
 2010 => "00010010",
 2011 => "00011000",
 2012 => "11011101",
 2013 => "01011001",
 2014 => "01110011",
 2015 => "01110010",
 2016 => "11110010",
 2017 => "01000001",
 2018 => "01100110",
 2019 => "00011111",
 2020 => "01111010",
 2021 => "01010101",
 2022 => "11100000",
 2023 => "01100100",
 2024 => "00001010",
 2025 => "01001000",
 2026 => "11110001",
 2027 => "10001110",
 2028 => "11011110",
 2029 => "00000010",
 2030 => "00011011",
 2031 => "10101100",
 2032 => "11000101",
 2033 => "11101101",
 2034 => "00011000",
 2035 => "00010111",
 2036 => "01100111",
 2037 => "01001111",
 2038 => "01010001",
 2039 => "01111001",
 2040 => "11001100",
 2041 => "11110000",
 2042 => "00101110",
 2043 => "01001110",
 2044 => "01111000",
 2045 => "00010010",
 2046 => "10111101",
 2047 => "01001111",
 2048 => "00011110",
 2049 => "11000100",
 2050 => "10001000",
 2051 => "00011111",
 2052 => "10111011",
 2053 => "00110101",
 2054 => "10101111",
 2055 => "10111100",
 2056 => "11110110",
 2057 => "00111111",
 2058 => "10001001",
 2059 => "01000100",
 2060 => "10000101",
 2061 => "00100010",
 2062 => "00010001",
 2063 => "01101010",
 2064 => "00110111",
 2065 => "00000011",
 2066 => "00111101",
 2067 => "10000110",
 2068 => "11001110",
 2069 => "01110001",
 2070 => "11101100",
 2071 => "00001000",
 2072 => "10010110",
 2073 => "11100010",
 2074 => "10011000",
 2075 => "01010001",
 2076 => "10011001",
 2077 => "01010010",
 2078 => "10100001",
 2079 => "00010101",
 2080 => "10110001",
 2081 => "00101101",
 2082 => "01010110",
 2083 => "10101111",
 2084 => "10101111",
 2085 => "00100001",
 2086 => "10111011",
 2087 => "01110111",
 2088 => "00111010",
 2089 => "11100111",
 2090 => "01011101",
 2091 => "00011000",
 2092 => "11000111",
 2093 => "00000011",
 2094 => "00101001",
 2095 => "11101111",
 2096 => "01100101",
 2097 => "10010101",
 2098 => "01111001",
 2099 => "00000010",
 2100 => "01100100",
 2101 => "01100010",
 2102 => "11000001",
 2103 => "10101110",
 2104 => "11100011",
 2105 => "10010111",
 2106 => "00111101",
 2107 => "00111101",
 2108 => "10001010",
 2109 => "10001110",
 2110 => "01000001",
 2111 => "00011010",
 2112 => "01110110",
 2113 => "01100111",
 2114 => "11010100",
 2115 => "01100001",
 2116 => "10001110",
 2117 => "00010110",
 2118 => "11111010",
 2119 => "10100101",
 2120 => "01101111",
 2121 => "01111000",
 2122 => "01100111",
 2123 => "11100100",
 2124 => "10110110",
 2125 => "01000111",
 2126 => "00101001",
 2127 => "10011010",
 2128 => "10000010",
 2129 => "00110111",
 2130 => "01000011",
 2131 => "11111101",
 2132 => "10001110",
 2133 => "10010100",
 2134 => "10001111",
 2135 => "00100100",
 2136 => "00110100",
 2137 => "00100000",
 2138 => "10011011",
 2139 => "10011101",
 2140 => "10110110",
 2141 => "11000011",
 2142 => "10101111",
 2143 => "01110100",
 2144 => "01011110",
 2145 => "00101001",
 2146 => "00011111",
 2147 => "10101111",
 2148 => "01001011",
 2149 => "00010001",
 2150 => "00001110",
 2151 => "10010100",
 2152 => "01111000",
 2153 => "10100110",
 2154 => "00010110",
 2155 => "11111110",
 2156 => "01011111",
 2157 => "00010100",
 2158 => "00111111",
 2159 => "01111011",
 2160 => "01010111",
 2161 => "10010001",
 2162 => "10100111",
 2163 => "01001111",
 2164 => "11100010",
 2165 => "11111100",
 2166 => "00011110",
 2167 => "11010000",
 2168 => "01001010",
 2169 => "01001100",
 2170 => "11001011",
 2171 => "00111111",
 2172 => "00100110",
 2173 => "11010000",
 2174 => "01011101",
 2175 => "00110000",
 2176 => "11101010",
 2177 => "01101011",
 2178 => "00011010",
 2179 => "11110010",
 2180 => "11100011",
 2181 => "10100101",
 2182 => "11001110",
 2183 => "01010111",
 2184 => "10111111",
 2185 => "10000010",
 2186 => "00000010",
 2187 => "10101101",
 2188 => "01000110",
 2189 => "11001011",
 2190 => "11111000",
 2191 => "01011011",
 2192 => "10111001",
 2193 => "11100100",
 2194 => "01111011",
 2195 => "11011011",
 2196 => "11100011",
 2197 => "01000101",
 2198 => "10111001",
 2199 => "10000100",
 2200 => "10111011",
 2201 => "01101011",
 2202 => "01010000",
 2203 => "01001011",
 2204 => "00111010",
 2205 => "00010001",
 2206 => "10100111",
 2207 => "11011001",
 2208 => "01111010",
 2209 => "10100111",
 2210 => "11001001",
 2211 => "10101001",
 2212 => "11100100",
 2213 => "11001101",
 2214 => "11011000",
 2215 => "00010011",
 2216 => "00111000",
 2217 => "10101101",
 2218 => "00011100",
 2219 => "00110011",
 2220 => "00010001",
 2221 => "01110101",
 2222 => "00111101",
 2223 => "01011010",
 2224 => "11110010",
 2225 => "01110000",
 2226 => "00000110",
 2227 => "10011011",
 2228 => "10100110",
 2229 => "11110110",
 2230 => "10100101",
 2231 => "00110111",
 2232 => "00011011",
 2233 => "11000111",
 2234 => "00100011",
 2235 => "10010001",
 2236 => "00100111",
 2237 => "01010110",
 2238 => "00100111",
 2239 => "01011010",
 2240 => "11001001",
 2241 => "11100011",
 2242 => "00100100",
 2243 => "01110010",
 2244 => "11110011",
 2245 => "10000110",
 2246 => "11100110",
 2247 => "01101100",
 2248 => "10110100",
 2249 => "11001010",
 2250 => "00001101",
 2251 => "00001010",
 2252 => "00111010",
 2253 => "10010010",
 2254 => "11110001",
 2255 => "10111011",
 2256 => "01100111",
 2257 => "11011010",
 2258 => "11010000",
 2259 => "01101001",
 2260 => "01001101",
 2261 => "10011101",
 2262 => "10100011",
 2263 => "10010001",
 2264 => "01110100",
 2265 => "00011001",
 2266 => "01001000",
 2267 => "01101111",
 2268 => "00110100",
 2269 => "11100010",
 2270 => "01011001",
 2271 => "11100010",
 2272 => "01100010",
 2273 => "10011101",
 2274 => "00110101",
 2275 => "01111100",
 2276 => "10000110",
 2277 => "10000000",
 2278 => "00100100",
 2279 => "01010001",
 2280 => "01111110",
 2281 => "10101011",
 2282 => "10000010",
 2283 => "01000010",
 2284 => "10001111",
 2285 => "01011010",
 2286 => "10100110",
 2287 => "10110000",
 2288 => "11010110",
 2289 => "11000000",
 2290 => "00101111",
 2291 => "00111000",
 2292 => "10100111",
 2293 => "10100110",
 2294 => "10101001",
 2295 => "01111100",
 2296 => "01111001",
 2297 => "00010000",
 2298 => "11000000",
 2299 => "01110011",
 2300 => "00110011",
 2301 => "11001100",
 2302 => "00001001",
 2303 => "11110011",
 2304 => "11111100",
 2305 => "01010110",
 2306 => "10100001",
 2307 => "01101010",
 2308 => "00011001",
 2309 => "10000100",
 2310 => "11001001",
 2311 => "11001011",
 2312 => "11010010",
 2313 => "00010101",
 2314 => "11110011",
 2315 => "10000010",
 2316 => "11010101",
 2317 => "01100001",
 2318 => "10100010",
 2319 => "11010100",
 2320 => "11011100",
 2321 => "00011111",
 2322 => "00001100",
 2323 => "00010100",
 2324 => "11111000",
 2325 => "11010110",
 2326 => "11101100",
 2327 => "11100001",
 2328 => "00111100",
 2329 => "00110111",
 2330 => "10011010",
 2331 => "11101110",
 2332 => "11011010",
 2333 => "10011100",
 2334 => "01111000",
 2335 => "01110000",
 2336 => "01100001",
 2337 => "10000011",
 2338 => "01011101",
 2339 => "01010101",
 2340 => "10001011",
 2341 => "01100111",
 2342 => "10101000",
 2343 => "11001001",
 2344 => "10000000",
 2345 => "11010000",
 2346 => "01101000",
 2347 => "11000001",
 2348 => "11011010",
 2349 => "01000110",
 2350 => "10101111",
 2351 => "00000001",
 2352 => "11111110",
 2353 => "10001100",
 2354 => "00010001",
 2355 => "00010010",
 2356 => "00010110",
 2357 => "00111101",
 2358 => "01101011",
 2359 => "01001010",
 2360 => "11110011",
 2361 => "10100101",
 2362 => "00101001",
 2363 => "10101011",
 2364 => "00110011",
 2365 => "11011001",
 2366 => "11001111",
 2367 => "01110011",
 2368 => "10101011",
 2369 => "01110000",
 2370 => "01010111",
 2371 => "10111010",
 2372 => "11000000",
 2373 => "01010101",
 2374 => "10001001",
 2375 => "00110110",
 2376 => "11010111",
 2377 => "11011000",
 2378 => "10111100",
 2379 => "10110000",
 2380 => "01010010",
 2381 => "00001010",
 2382 => "10011111",
 2383 => "11101011",
 2384 => "11101010",
 2385 => "01111100",
 2386 => "01110110",
 2387 => "00000101",
 2388 => "11111011",
 2389 => "01010111",
 2390 => "00110011",
 2391 => "10110000",
 2392 => "00100001",
 2393 => "11101110",
 2394 => "00111011",
 2395 => "10001011",
 2396 => "00111111",
 2397 => "11111000",
 2398 => "10110011",
 2399 => "10110111",
 2400 => "10101001",
 2401 => "11101100",
 2402 => "10000001",
 2403 => "10111001",
 2404 => "11011010",
 2405 => "00110000",
 2406 => "11100100",
 2407 => "01010100",
 2408 => "10111110",
 2409 => "10010000",
 2410 => "11111100",
 2411 => "00000001",
 2412 => "00100010",
 2413 => "00111100",
 2414 => "10100001",
 2415 => "01000111",
 2416 => "10011111",
 2417 => "10111010",
 2418 => "11000011",
 2419 => "01011110",
 2420 => "11011101",
 2421 => "00011110",
 2422 => "00011100",
 2423 => "11011001",
 2424 => "10111111",
 2425 => "10100011",
 2426 => "11100100",
 2427 => "10101010",
 2428 => "11101011",
 2429 => "10010001",
 2430 => "10100011",
 2431 => "11101011",
 2432 => "10101011",
 2433 => "01110110",
 2434 => "00100010",
 2435 => "10001000",
 2436 => "10010010",
 2437 => "10110111",
 2438 => "10001010",
 2439 => "11011100",
 2440 => "10110000",
 2441 => "00010111",
 2442 => "00110101",
 2443 => "01001011",
 2444 => "11101010",
 2445 => "01001101",
 2446 => "11101001",
 2447 => "00111110",
 2448 => "10101010",
 2449 => "01001000",
 2450 => "00101101",
 2451 => "00011001",
 2452 => "10001010",
 2453 => "10111011",
 2454 => "01001100",
 2455 => "01000000",
 2456 => "11101100",
 2457 => "01110110",
 2458 => "01100101",
 2459 => "11000010",
 2460 => "01100001",
 2461 => "11111111",
 2462 => "10100100",
 2463 => "01101000",
 2464 => "00011010",
 2465 => "10111101",
 2466 => "10101111",
 2467 => "00100000",
 2468 => "11010111",
 2469 => "11101011",
 2470 => "01111001",
 2471 => "11001110",
 2472 => "11001101",
 2473 => "00100010",
 2474 => "10001010",
 2475 => "01101000",
 2476 => "01111111",
 2477 => "01111010",
 2478 => "01110000",
 2479 => "00001110",
 2480 => "11010110",
 2481 => "10000110",
 2482 => "01100100",
 2483 => "00111101",
 2484 => "01011000",
 2485 => "01001101",
 2486 => "11110010",
 2487 => "00110111",
 2488 => "01000001",
 2489 => "01100001",
 2490 => "11110111",
 2491 => "01100101",
 2492 => "00101000",
 2493 => "11111011",
 2494 => "11111111",
 2495 => "00101010",
 2496 => "00100000",
 2497 => "10101010",
 2498 => "01000101",
 2499 => "10001000",
 2500 => "11100110",
 2501 => "10111110",
 2502 => "00011101",
 2503 => "01110011",
 2504 => "10000010",
 2505 => "10110111",
 2506 => "11110111",
 2507 => "01101101",
 2508 => "00100000",
 2509 => "11100011",
 2510 => "10000101",
 2511 => "11100001",
 2512 => "11010001",
 2513 => "10010010",
 2514 => "00010100",
 2515 => "00111011",
 2516 => "00100100",
 2517 => "11001111",
 2518 => "00110011",
 2519 => "01011001",
 2520 => "11101100",
 2521 => "11101001",
 2522 => "10110100",
 2523 => "10110101",
 2524 => "00001101",
 2525 => "10111110",
 2526 => "10001001",
 2527 => "00000010",
 2528 => "10110001",
 2529 => "10101010",
 2530 => "10011111",
 2531 => "10010110",
 2532 => "11110011",
 2533 => "01101011",
 2534 => "01011000",
 2535 => "01110101",
 2536 => "01101011",
 2537 => "11101001",
 2538 => "00110100",
 2539 => "00011010",
 2540 => "01110011",
 2541 => "01011110",
 2542 => "10000000",
 2543 => "10111101",
 2544 => "10001011",
 2545 => "00000000",
 2546 => "11001111",
 2547 => "00101010",
 2548 => "01110100",
 2549 => "01110111",
 2550 => "00001110",
 2551 => "11011111",
 2552 => "00010001",
 2553 => "10100110",
 2554 => "00000011",
 2555 => "10011101",
 2556 => "10101000",
 2557 => "01001100",
 2558 => "10100011",
 2559 => "00010010",
 2560 => "11011110",
 2561 => "11100110",
 2562 => "11000010",
 2563 => "11111010",
 2564 => "11111101",
 2565 => "10111111",
 2566 => "01111110",
 2567 => "00000111",
 2568 => "01110011",
 2569 => "10000000",
 2570 => "11110101",
 2571 => "11100111",
 2572 => "10000000",
 2573 => "00110111",
 2574 => "10111000",
 2575 => "00100111",
 2576 => "01100100",
 2577 => "11111110",
 2578 => "01011000",
 2579 => "10101100",
 2580 => "00110110",
 2581 => "00001001",
 2582 => "01010010",
 2583 => "01110011",
 2584 => "01110111",
 2585 => "00110100",
 2586 => "11000001",
 2587 => "10111111",
 2588 => "10001110",
 2589 => "00000110",
 2590 => "01100110",
 2591 => "01000001",
 2592 => "10010111",
 2593 => "11110001",
 2594 => "00000011",
 2595 => "00101011",
 2596 => "01011010",
 2597 => "00000110",
 2598 => "00110001",
 2599 => "11000010",
 2600 => "00110111",
 2601 => "01000010",
 2602 => "00010011",
 2603 => "11100111",
 2604 => "01111010",
 2605 => "10000011",
 2606 => "00100100",
 2607 => "10001100",
 2608 => "11001111",
 2609 => "01001100",
 2610 => "00000101",
 2611 => "10000001",
 2612 => "10101101",
 2613 => "11010100",
 2614 => "00111101",
 2615 => "10110001",
 2616 => "10011111",
 2617 => "01110111",
 2618 => "10001101",
 2619 => "11100001",
 2620 => "01110110",
 2621 => "00111000",
 2622 => "10100111",
 2623 => "10110100",
 2624 => "10000110",
 2625 => "01001001",
 2626 => "11100100",
 2627 => "11001111",
 2628 => "00001011",
 2629 => "10110001",
 2630 => "10100100",
 2631 => "11111111",
 2632 => "01010000",
 2633 => "10110101",
 2634 => "10110011",
 2635 => "10011101",
 2636 => "01010111",
 2637 => "01110111",
 2638 => "10010010",
 2639 => "01000101",
 2640 => "00000000",
 2641 => "10010000",
 2642 => "11100111",
 2643 => "01100111",
 2644 => "01110101",
 2645 => "00000001",
 2646 => "11011010",
 2647 => "11001100",
 2648 => "11001111",
 2649 => "01101010",
 2650 => "11101110",
 2651 => "11010010",
 2652 => "10100000",
 2653 => "01100000",
 2654 => "00100011",
 2655 => "11001110",
 2656 => "00101010",
 2657 => "11000010",
 2658 => "11010011",
 2659 => "10011011",
 2660 => "00001101",
 2661 => "00000100",
 2662 => "10100001",
 2663 => "01111000",
 2664 => "11010000",
 2665 => "00111100",
 2666 => "01100010",
 2667 => "10001110",
 2668 => "11100010",
 2669 => "01001100",
 2670 => "00010001",
 2671 => "11000000",
 2672 => "10101110",
 2673 => "10001000",
 2674 => "10111010",
 2675 => "10000101",
 2676 => "01010100",
 2677 => "11101100",
 2678 => "11011000",
 2679 => "01110100",
 2680 => "10111101",
 2681 => "10010101",
 2682 => "00101111",
 2683 => "01101111",
 2684 => "00011010",
 2685 => "11101101",
 2686 => "11000100",
 2687 => "11110001",
 2688 => "11111101",
 2689 => "10100001",
 2690 => "00100000",
 2691 => "00101000",
 2692 => "11100000",
 2693 => "11100001",
 2694 => "10000111",
 2695 => "00000011",
 2696 => "10100001",
 2697 => "00000001",
 2698 => "00111011",
 2699 => "01101110",
 2700 => "10010001",
 2701 => "10011100",
 2702 => "11111101",
 2703 => "10100001",
 2704 => "00011000",
 2705 => "01001010",
 2706 => "01010010",
 2707 => "00100001",
 2708 => "00010001",
 2709 => "11100010",
 2710 => "11101110",
 2711 => "01111111",
 2712 => "00010011",
 2713 => "11000101",
 2714 => "00110101",
 2715 => "10111100",
 2716 => "11011101",
 2717 => "10100000",
 2718 => "10001111",
 2719 => "00111000",
 2720 => "01011111",
 2721 => "00110111",
 2722 => "01001111",
 2723 => "00001110",
 2724 => "00101111",
 2725 => "01110100",
 2726 => "00110001",
 2727 => "10010111",
 2728 => "00110000",
 2729 => "11100101",
 2730 => "01011000",
 2731 => "10101010",
 2732 => "01001110",
 2733 => "11001100",
 2734 => "00011001",
 2735 => "00111101",
 2736 => "00001000",
 2737 => "00011011",
 2738 => "10001101",
 2739 => "10001110",
 2740 => "00101000",
 2741 => "11111010",
 2742 => "01011011",
 2743 => "11000111",
 2744 => "10100011",
 2745 => "00100101",
 2746 => "10101000",
 2747 => "00111101",
 2748 => "11101111",
 2749 => "10110001",
 2750 => "01010100",
 2751 => "11001100",
 2752 => "11111010",
 2753 => "01100100",
 2754 => "00000101",
 2755 => "10001110",
 2756 => "00100101",
 2757 => "00000001",
 2758 => "01111000",
 2759 => "10100101",
 2760 => "00110100",
 2761 => "00100110",
 2762 => "10100000",
 2763 => "10111111",
 2764 => "00001010",
 2765 => "01011101",
 2766 => "10001100",
 2767 => "10100110",
 2768 => "00001010",
 2769 => "11111011",
 2770 => "10000110",
 2771 => "00011000",
 2772 => "01000101",
 2773 => "10110011",
 2774 => "10011100",
 2775 => "11010100",
 2776 => "10100011",
 2777 => "01001111",
 2778 => "11001011",
 2779 => "11011000",
 2780 => "00101110",
 2781 => "10110010",
 2782 => "11100001",
 2783 => "10100011",
 2784 => "01100101",
 2785 => "00100010",
 2786 => "10001010",
 2787 => "10101111",
 2788 => "10010100",
 2789 => "00011011",
 2790 => "00000111",
 2791 => "11101110",
 2792 => "10111011",
 2793 => "11001101",
 2794 => "00101110",
 2795 => "11100001",
 2796 => "11100101",
 2797 => "01011110",
 2798 => "00000011",
 2799 => "11000001",
 2800 => "11010111",
 2801 => "11111001",
 2802 => "11011110",
 2803 => "11010000",
 2804 => "10010011",
 2805 => "00100100",
 2806 => "01010101",
 2807 => "01111011",
 2808 => "11011001",
 2809 => "11101001",
 2810 => "00100110",
 2811 => "11100011",
 2812 => "10000111",
 2813 => "10110011",
 2814 => "00010110",
 2815 => "11100011",
 2816 => "10110100",
 2817 => "01010011",
 2818 => "11111101",
 2819 => "01100011",
 2820 => "01111010",
 2821 => "10110000",
 2822 => "11100101",
 2823 => "11100011",
 2824 => "10001110",
 2825 => "00000011",
 2826 => "11111110",
 2827 => "01100001",
 2828 => "01010011",
 2829 => "11000010",
 2830 => "01010111",
 2831 => "10111001",
 2832 => "10100101",
 2833 => "11010010",
 2834 => "00111110",
 2835 => "01000001",
 2836 => "11010001",
 2837 => "00110010",
 2838 => "01111001",
 2839 => "11011001",
 2840 => "00000011",
 2841 => "00100000",
 2842 => "01101001",
 2843 => "11110101",
 2844 => "10001010",
 2845 => "00010000",
 2846 => "11010101",
 2847 => "01110000",
 2848 => "10101110",
 2849 => "00000110",
 2850 => "01000100",
 2851 => "00010101",
 2852 => "01010010",
 2853 => "01011000",
 2854 => "10111110",
 2855 => "01110000",
 2856 => "00001101",
 2857 => "11011111",
 2858 => "11011111",
 2859 => "10000101",
 2860 => "01111101",
 2861 => "11001101",
 2862 => "11010001",
 2863 => "11110101",
 2864 => "01101001",
 2865 => "11110101",
 2866 => "01001110",
 2867 => "10001111",
 2868 => "00010110",
 2869 => "11110111",
 2870 => "10001010",
 2871 => "11000101",
 2872 => "10111001",
 2873 => "01000111",
 2874 => "00111011",
 2875 => "01110000",
 2876 => "11011000",
 2877 => "11000011",
 2878 => "10010010",
 2879 => "11010010",
 2880 => "10010110",
 2881 => "10001001",
 2882 => "00100100",
 2883 => "00001101",
 2884 => "11100111",
 2885 => "01100111",
 2886 => "01111110",
 2887 => "00100111",
 2888 => "01001001",
 2889 => "00100111",
 2890 => "11010101",
 2891 => "00011101",
 2892 => "01011000",
 2893 => "00001011",
 2894 => "11000111",
 2895 => "11101110",
 2896 => "11000010",
 2897 => "01100011",
 2898 => "11001011",
 2899 => "10101110",
 2900 => "11010111",
 2901 => "00000111",
 2902 => "00011101",
 2903 => "10000110",
 2904 => "00001100",
 2905 => "00100101",
 2906 => "11101000",
 2907 => "10000111",
 2908 => "11111010",
 2909 => "01011000",
 2910 => "11110010",
 2911 => "11001101",
 2912 => "11001101",
 2913 => "00010001",
 2914 => "00000011",
 2915 => "11110110",
 2916 => "00001101",
 2917 => "01111111",
 2918 => "01001110",
 2919 => "10110001",
 2920 => "01010101",
 2921 => "00000111",
 2922 => "10000001",
 2923 => "01111010",
 2924 => "11010000",
 2925 => "00101110",
 2926 => "01111110",
 2927 => "00100111",
 2928 => "10111000",
 2929 => "10101110",
 2930 => "11110101",
 2931 => "10011010",
 2932 => "10011101",
 2933 => "00111000",
 2934 => "00001001",
 2935 => "01000000",
 2936 => "10001100",
 2937 => "11111111",
 2938 => "01111100",
 2939 => "00111111",
 2940 => "10100110",
 2941 => "01111000",
 2942 => "01100110",
 2943 => "01101010",
 2944 => "10111011",
 2945 => "00101001",
 2946 => "01110101",
 2947 => "01100111",
 2948 => "00111010",
 2949 => "11000000",
 2950 => "00001001",
 2951 => "10101000",
 2952 => "01100001",
 2953 => "00011100",
 2954 => "10011010",
 2955 => "11111101",
 2956 => "10100000",
 2957 => "00101010",
 2958 => "01011001",
 2959 => "10110000",
 2960 => "00010011",
 2961 => "10000100",
 2962 => "11010110",
 2963 => "01001110",
 2964 => "01100011",
 2965 => "10011010",
 2966 => "11000101",
 2967 => "01000000",
 2968 => "10000111",
 2969 => "01010100",
 2970 => "00100100",
 2971 => "10011011",
 2972 => "01010111",
 2973 => "11110111",
 2974 => "10101100",
 2975 => "00100011",
 2976 => "01001001",
 2977 => "00010001",
 2978 => "01110001",
 2979 => "01011010",
 2980 => "10100110",
 2981 => "10010100",
 2982 => "11101000",
 2983 => "00000100",
 2984 => "00000110",
 2985 => "00101001",
 2986 => "10111011",
 2987 => "10100110",
 2988 => "11100100",
 2989 => "01001100",
 2990 => "01011110",
 2991 => "11011011",
 2992 => "11001001",
 2993 => "10001010",
 2994 => "01111011",
 2995 => "11111001",
 2996 => "01011001",
 2997 => "11000011",
 2998 => "11111100",
 2999 => "01000100",
 3000 => "01101011",
 3001 => "10001110",
 3002 => "11001000",
 3003 => "10000101",
 3004 => "10111110",
 3005 => "10100010",
 3006 => "01101110",
 3007 => "11001000",
 3008 => "10110001",
 3009 => "10011011",
 3010 => "00010011",
 3011 => "10010101",
 3012 => "00101100",
 3013 => "11111011",
 3014 => "11001100",
 3015 => "11100100",
 3016 => "01101010",
 3017 => "10100101",
 3018 => "11111001",
 3019 => "11011100",
 3020 => "01010101",
 3021 => "00100000",
 3022 => "11111000",
 3023 => "00101111",
 3024 => "10110101",
 3025 => "10011001",
 3026 => "10110000",
 3027 => "10101011",
 3028 => "00101110",
 3029 => "10111001",
 3030 => "00100000",
 3031 => "01101101",
 3032 => "00011000",
 3033 => "11010101",
 3034 => "01100001",
 3035 => "00010010",
 3036 => "01100110",
 3037 => "10100001",
 3038 => "10110011",
 3039 => "11000111",
 3040 => "01110000",
 3041 => "11011110",
 3042 => "01010111",
 3043 => "00000100",
 3044 => "10011010",
 3045 => "10010101",
 3046 => "10111011",
 3047 => "01111011",
 3048 => "00010010",
 3049 => "00001100",
 3050 => "00100110",
 3051 => "01000110",
 3052 => "00110111",
 3053 => "10001111",
 3054 => "11110111",
 3055 => "10101100",
 3056 => "10000110",
 3057 => "11010110",
 3058 => "10101001",
 3059 => "00011110",
 3060 => "11111010",
 3061 => "01101011",
 3062 => "01101100",
 3063 => "01101001",
 3064 => "01010101",
 3065 => "11010101",
 3066 => "11111110",
 3067 => "00000001",
 3068 => "01010100",
 3069 => "11011101",
 3070 => "01100001",
 3071 => "10000000",
 3072 => "11111110",
 3073 => "11110111",
 3074 => "10000101",
 3075 => "10111000",
 3076 => "10000001",
 3077 => "01010011",
 3078 => "11101001",
 3079 => "00101010",
 3080 => "10110110",
 3081 => "00011101",
 3082 => "11000010",
 3083 => "10010010",
 3084 => "11011101",
 3085 => "01001000",
 3086 => "11111100",
 3087 => "11000011",
 3088 => "00101000",
 3089 => "00111010",
 3090 => "00000000",
 3091 => "11111011",
 3092 => "01110010",
 3093 => "01111100",
 3094 => "01101010",
 3095 => "01010101",
 3096 => "10101111",
 3097 => "11111111",
 3098 => "00111101",
 3099 => "10001001",
 3100 => "01001010",
 3101 => "10000100",
 3102 => "01001111",
 3103 => "11000001",
 3104 => "01010011",
 3105 => "10110110",
 3106 => "10001111",
 3107 => "00011000",
 3108 => "00000000",
 3109 => "01100100",
 3110 => "10110111",
 3111 => "01001101",
 3112 => "01100010",
 3113 => "11111000",
 3114 => "10101111",
 3115 => "01000001",
 3116 => "10101110",
 3117 => "10001111",
 3118 => "10010110",
 3119 => "11000011",
 3120 => "11011110",
 3121 => "11011100",
 3122 => "01100101",
 3123 => "01000101",
 3124 => "10010100",
 3125 => "01101000",
 3126 => "01111001",
 3127 => "01000000",
 3128 => "11001011",
 3129 => "11100101",
 3130 => "11101110",
 3131 => "11011110",
 3132 => "00010001",
 3133 => "01110001",
 3134 => "01110101",
 3135 => "00001000",
 3136 => "01001110",
 3137 => "01001001",
 3138 => "00000000",
 3139 => "00000001",
 3140 => "10110100",
 3141 => "00111100",
 3142 => "00011010",
 3143 => "01101011",
 3144 => "10100101",
 3145 => "11001010",
 3146 => "11000010",
 3147 => "00111011",
 3148 => "11000110",
 3149 => "01101111",
 3150 => "10011110",
 3151 => "00000001",
 3152 => "00100000",
 3153 => "10111101",
 3154 => "00001011",
 3155 => "01101000",
 3156 => "10101111",
 3157 => "01000010",
 3158 => "10100111",
 3159 => "01000111",
 3160 => "11010110",
 3161 => "01011111",
 3162 => "11011000",
 3163 => "11001100",
 3164 => "10110111",
 3165 => "10010111",
 3166 => "01110100",
 3167 => "10110111",
 3168 => "00000010",
 3169 => "01100000",
 3170 => "00111011",
 3171 => "00000001",
 3172 => "00100111",
 3173 => "11100111",
 3174 => "10010110",
 3175 => "00101110",
 3176 => "11001110",
 3177 => "11110011",
 3178 => "01110101",
 3179 => "00110100",
 3180 => "10010101",
 3181 => "01100011",
 3182 => "01010011",
 3183 => "00001010",
 3184 => "10100010",
 3185 => "00000011",
 3186 => "10100000",
 3187 => "01000011",
 3188 => "01110010",
 3189 => "11110100",
 3190 => "00011000",
 3191 => "10010011",
 3192 => "10001000",
 3193 => "01000001",
 3194 => "10001101",
 3195 => "11010011",
 3196 => "10110010",
 3197 => "01010111",
 3198 => "10100010",
 3199 => "10100110",
 3200 => "10100101",
 3201 => "01011011",
 3202 => "10011101",
 3203 => "01101110",
 3204 => "00111100",
 3205 => "11010100",
 3206 => "11000011",
 3207 => "11111011",
 3208 => "00111110",
 3209 => "01001110",
 3210 => "10011000",
 3211 => "01010000",
 3212 => "10101110",
 3213 => "00011100",
 3214 => "01100101",
 3215 => "00000111",
 3216 => "01011110",
 3217 => "01110000",
 3218 => "01110011",
 3219 => "10001111",
 3220 => "00010100",
 3221 => "01100000",
 3222 => "00011000",
 3223 => "01101111",
 3224 => "11000100",
 3225 => "00100110",
 3226 => "01011101",
 3227 => "11000010",
 3228 => "10101000",
 3229 => "01110101",
 3230 => "01000101",
 3231 => "11111100",
 3232 => "10010111",
 3233 => "11100000",
 3234 => "10011011",
 3235 => "01010011",
 3236 => "10111000",
 3237 => "01011001",
 3238 => "10011010",
 3239 => "11000000",
 3240 => "00001110",
 3241 => "10111000",
 3242 => "01011000",
 3243 => "11011110",
 3244 => "01001000",
 3245 => "10101110",
 3246 => "10110000",
 3247 => "11110100",
 3248 => "00101110",
 3249 => "10111101",
 3250 => "11110110",
 3251 => "10111010",
 3252 => "11010000",
 3253 => "00010011",
 3254 => "01000110",
 3255 => "00011001",
 3256 => "11011111",
 3257 => "00100111",
 3258 => "01101110",
 3259 => "10101000",
 3260 => "00010110",
 3261 => "10010101",
 3262 => "00000001",
 3263 => "01001110",
 3264 => "00011010",
 3265 => "01011011",
 3266 => "11011011",
 3267 => "10111100",
 3268 => "10101011",
 3269 => "11000101",
 3270 => "11111110",
 3271 => "10101011",
 3272 => "10000111",
 3273 => "10010011",
 3274 => "01100110",
 3275 => "11101110",
 3276 => "00100111",
 3277 => "10011101",
 3278 => "01010101",
 3279 => "01111100",
 3280 => "11001110",
 3281 => "01011000",
 3282 => "01101000",
 3283 => "10110100",
 3284 => "01010000",
 3285 => "00011101",
 3286 => "00000110",
 3287 => "10110110",
 3288 => "01100100",
 3289 => "11001010",
 3290 => "10111000",
 3291 => "11010011",
 3292 => "10111100",
 3293 => "01110101",
 3294 => "10111110",
 3295 => "01110110",
 3296 => "11001001",
 3297 => "11111111",
 3298 => "11101000",
 3299 => "01011100",
 3300 => "01100101",
 3301 => "11111001",
 3302 => "11010110",
 3303 => "10010011",
 3304 => "01100001",
 3305 => "01011011",
 3306 => "10001011",
 3307 => "11101011",
 3308 => "00111011",
 3309 => "11111100",
 3310 => "11110100",
 3311 => "11111111",
 3312 => "01101110",
 3313 => "10100011",
 3314 => "00000111",
 3315 => "11001101",
 3316 => "01110011",
 3317 => "01100111",
 3318 => "01010100",
 3319 => "00000000",
 3320 => "00100100",
 3321 => "10101010",
 3322 => "01100011",
 3323 => "11110100",
 3324 => "01111001",
 3325 => "10000010",
 3326 => "10010101",
 3327 => "10101111",
 3328 => "10000001",
 3329 => "11100011",
 3330 => "11010110",
 3331 => "10010100",
 3332 => "01100100",
 3333 => "11110000",
 3334 => "11100011",
 3335 => "00001110",
 3336 => "11100001",
 3337 => "10001111",
 3338 => "11110101",
 3339 => "11100110",
 3340 => "10011111",
 3341 => "01011010",
 3342 => "01010101",
 3343 => "10100100",
 3344 => "10110000",
 3345 => "11111000",
 3346 => "00011001",
 3347 => "01001000",
 3348 => "10100101",
 3349 => "00001110",
 3350 => "01100010",
 3351 => "00011100",
 3352 => "11000000",
 3353 => "10010110",
 3354 => "00010111",
 3355 => "01100101",
 3356 => "00001101",
 3357 => "10100000",
 3358 => "01011000",
 3359 => "10011001",
 3360 => "00001001",
 3361 => "00101101",
 3362 => "10000010",
 3363 => "10100100",
 3364 => "10100001",
 3365 => "10110000",
 3366 => "00100110",
 3367 => "01011010",
 3368 => "11100011",
 3369 => "00101001",
 3370 => "01000010",
 3371 => "10111000",
 3372 => "00101110",
 3373 => "00100011",
 3374 => "00100010",
 3375 => "00000101",
 3376 => "10001000",
 3377 => "01011110",
 3378 => "00010111",
 3379 => "00000011",
 3380 => "01111010",
 3381 => "01101110",
 3382 => "00001010",
 3383 => "11000000",
 3384 => "01110110",
 3385 => "01101101",
 3386 => "00101010",
 3387 => "10101100",
 3388 => "10000101",
 3389 => "00010011",
 3390 => "00100110",
 3391 => "00100001",
 3392 => "00111011",
 3393 => "01001000",
 3394 => "01111001",
 3395 => "11000000",
 3396 => "01110101",
 3397 => "01011111",
 3398 => "00010100",
 3399 => "10110011",
 3400 => "00011101",
 3401 => "10010101",
 3402 => "11001000",
 3403 => "11000011",
 3404 => "00111111",
 3405 => "10110011",
 3406 => "11001100",
 3407 => "10111010",
 3408 => "01001001",
 3409 => "11101110",
 3410 => "10110000",
 3411 => "10001000",
 3412 => "01001011",
 3413 => "11011010",
 3414 => "01100001",
 3415 => "11011111",
 3416 => "10110111",
 3417 => "11011110",
 3418 => "00100110",
 3419 => "10000101",
 3420 => "01000101",
 3421 => "10010100",
 3422 => "00101010",
 3423 => "11000011",
 3424 => "00111110",
 3425 => "10101101",
 3426 => "10010110",
 3427 => "00000111",
 3428 => "10000000",
 3429 => "01100111",
 3430 => "01000010",
 3431 => "11011001",
 3432 => "00001011",
 3433 => "01000000",
 3434 => "11011101",
 3435 => "11111010",
 3436 => "00110001",
 3437 => "00001111",
 3438 => "01010111",
 3439 => "01001001",
 3440 => "11101110",
 3441 => "10101011",
 3442 => "01011101",
 3443 => "00111001",
 3444 => "00101010",
 3445 => "10010100",
 3446 => "01101000",
 3447 => "00000000",
 3448 => "01101010",
 3449 => "01110111",
 3450 => "00000110",
 3451 => "11001010",
 3452 => "11010100",
 3453 => "10101001",
 3454 => "10011110",
 3455 => "01010000",
 3456 => "00110101",
 3457 => "11010010",
 3458 => "01000101",
 3459 => "10000100",
 3460 => "11111110",
 3461 => "01011100",
 3462 => "11010101",
 3463 => "10110001",
 3464 => "11101000",
 3465 => "11011100",
 3466 => "10100001",
 3467 => "10110011",
 3468 => "00001101",
 3469 => "10101111",
 3470 => "00100011",
 3471 => "00000001",
 3472 => "00011100",
 3473 => "00111011",
 3474 => "01111111",
 3475 => "11011110",
 3476 => "10100011",
 3477 => "11100001",
 3478 => "01110001",
 3479 => "01100111",
 3480 => "11010011",
 3481 => "00001000",
 3482 => "01101111",
 3483 => "10101101",
 3484 => "10100100",
 3485 => "01011101",
 3486 => "11101100",
 3487 => "01101101",
 3488 => "11110001",
 3489 => "11101110",
 3490 => "00111000",
 3491 => "10100111",
 3492 => "11110111",
 3493 => "01001010",
 3494 => "11011110",
 3495 => "11001001",
 3496 => "00000111",
 3497 => "11100010",
 3498 => "11010010",
 3499 => "00000101",
 3500 => "00011011",
 3501 => "00110101",
 3502 => "00111101",
 3503 => "10110001",
 3504 => "01100101",
 3505 => "01100010",
 3506 => "00111101",
 3507 => "00001101",
 3508 => "11001000",
 3509 => "11111011",
 3510 => "00011100",
 3511 => "10111010",
 3512 => "10101010",
 3513 => "01000001",
 3514 => "11100011",
 3515 => "00011100",
 3516 => "10001101",
 3517 => "01100111",
 3518 => "00001110",
 3519 => "00110011",
 3520 => "01111010",
 3521 => "10010110",
 3522 => "00101001",
 3523 => "01000110",
 3524 => "11010110",
 3525 => "11110010",
 3526 => "01110011",
 3527 => "01001101",
 3528 => "00111001",
 3529 => "01100110",
 3530 => "10010001",
 3531 => "10011000",
 3532 => "00010010",
 3533 => "01111010",
 3534 => "00001001",
 3535 => "11101101",
 3536 => "10010111",
 3537 => "01101010",
 3538 => "10100110",
 3539 => "01010011",
 3540 => "10000000",
 3541 => "00010111",
 3542 => "01010001",
 3543 => "00111011",
 3544 => "11110001",
 3545 => "01110011",
 3546 => "01111010",
 3547 => "11110010",
 3548 => "01101111",
 3549 => "11000111",
 3550 => "10111110",
 3551 => "10111001",
 3552 => "10011101",
 3553 => "11000010",
 3554 => "10011000",
 3555 => "00110010",
 3556 => "11001101",
 3557 => "11101110",
 3558 => "00000000",
 3559 => "00010101",
 3560 => "11111001",
 3561 => "00010101",
 3562 => "00110010",
 3563 => "11111010",
 3564 => "01011010",
 3565 => "01111111",
 3566 => "01010100",
 3567 => "01101000",
 3568 => "10001000",
 3569 => "01000111",
 3570 => "00010010",
 3571 => "11010000",
 3572 => "10100000",
 3573 => "01101101",
 3574 => "01100011",
 3575 => "11100101",
 3576 => "01000000",
 3577 => "11101111",
 3578 => "00001100",
 3579 => "11001000",
 3580 => "10000000",
 3581 => "00100101",
 3582 => "01111000",
 3583 => "10101000",
 3584 => "11001110",
 3585 => "10111011",
 3586 => "10110011",
 3587 => "11000100",
 3588 => "11101110",
 3589 => "11010000",
 3590 => "00101101",
 3591 => "10110000",
 3592 => "11101010",
 3593 => "01101101",
 3594 => "10100111",
 3595 => "10101000",
 3596 => "00000001",
 3597 => "01101010",
 3598 => "00000011",
 3599 => "01000110",
 3600 => "11011111",
 3601 => "10101101",
 3602 => "10000111",
 3603 => "00110001",
 3604 => "01110101",
 3605 => "11101110",
 3606 => "01011000",
 3607 => "10011011",
 3608 => "00011001",
 3609 => "01010100",
 3610 => "01000100",
 3611 => "10000110",
 3612 => "00100110",
 3613 => "10001110",
 3614 => "11111010",
 3615 => "11010101",
 3616 => "10001101",
 3617 => "11001111",
 3618 => "01100001",
 3619 => "10110101",
 3620 => "11111110",
 3621 => "10110001",
 3622 => "11010110",
 3623 => "00001111",
 3624 => "01101110",
 3625 => "10011011",
 3626 => "01101111",
 3627 => "11000000",
 3628 => "11000000",
 3629 => "01000001",
 3630 => "00100011",
 3631 => "10001010",
 3632 => "01000101",
 3633 => "11101110",
 3634 => "10111011",
 3635 => "00011100",
 3636 => "11111011",
 3637 => "10111011",
 3638 => "01001111",
 3639 => "11101101",
 3640 => "01100101",
 3641 => "00110011",
 3642 => "00001001",
 3643 => "01101010",
 3644 => "10000111",
 3645 => "10101010",
 3646 => "01010000",
 3647 => "10110111",
 3648 => "00101011",
 3649 => "01100010",
 3650 => "01111110",
 3651 => "00001110",
 3652 => "00110111",
 3653 => "01110101",
 3654 => "11101011",
 3655 => "00111010",
 3656 => "11001110",
 3657 => "01101100",
 3658 => "11001110",
 3659 => "10001000",
 3660 => "01000001",
 3661 => "11001001",
 3662 => "11111000",
 3663 => "11111011",
 3664 => "01111111",
 3665 => "00011110",
 3666 => "01110011",
 3667 => "00110011",
 3668 => "00011111",
 3669 => "01101100",
 3670 => "01100000",
 3671 => "10000001",
 3672 => "01011001",
 3673 => "01010100",
 3674 => "10011110",
 3675 => "11101111",
 3676 => "11010110",
 3677 => "01101001",
 3678 => "00111011",
 3679 => "01001011",
 3680 => "01101100",
 3681 => "00001111",
 3682 => "00010001",
 3683 => "11000000",
 3684 => "11001011",
 3685 => "00011000",
 3686 => "10100011",
 3687 => "00010010",
 3688 => "00011110",
 3689 => "00011110",
 3690 => "11101011",
 3691 => "01010000",
 3692 => "00000010",
 3693 => "01010011",
 3694 => "10100111",
 3695 => "11000110",
 3696 => "10011111",
 3697 => "01100011",
 3698 => "00110111",
 3699 => "10110100",
 3700 => "00000010",
 3701 => "01011011",
 3702 => "10111110",
 3703 => "10010001",
 3704 => "10000110",
 3705 => "01110100",
 3706 => "00011001",
 3707 => "00000001",
 3708 => "01011011",
 3709 => "10110110",
 3710 => "10000110",
 3711 => "01001110",
 3712 => "00000001",
 3713 => "01010001",
 3714 => "00001011",
 3715 => "00011110",
 3716 => "11101101",
 3717 => "11011110",
 3718 => "11101101",
 3719 => "00101100",
 3720 => "10110011",
 3721 => "10011110",
 3722 => "01011010",
 3723 => "01101001",
 3724 => "10110001",
 3725 => "00000101",
 3726 => "11001101",
 3727 => "00000110",
 3728 => "10100101",
 3729 => "10010000",
 3730 => "11011100",
 3731 => "10011101",
 3732 => "10110000",
 3733 => "11001101",
 3734 => "11010111",
 3735 => "00000111",
 3736 => "00110011",
 3737 => "10100111",
 3738 => "11111100",
 3739 => "01110001",
 3740 => "01011110",
 3741 => "00010011",
 3742 => "10111100",
 3743 => "11000110",
 3744 => "10100100",
 3745 => "00011100",
 3746 => "11000100",
 3747 => "00000100",
 3748 => "01101010",
 3749 => "00010110",
 3750 => "11100000",
 3751 => "11110001",
 3752 => "00001010",
 3753 => "11100111",
 3754 => "00011110",
 3755 => "00101011",
 3756 => "01010010",
 3757 => "11010001",
 3758 => "00010000",
 3759 => "01010001",
 3760 => "10100000",
 3761 => "00000001",
 3762 => "10100001",
 3763 => "10110010",
 3764 => "01111011",
 3765 => "01110000",
 3766 => "11101100",
 3767 => "01101011",
 3768 => "11101001",
 3769 => "10101000",
 3770 => "01010100",
 3771 => "00010010",
 3772 => "00100000",
 3773 => "00001111",
 3774 => "00110110",
 3775 => "11010000",
 3776 => "00100110",
 3777 => "00010001",
 3778 => "00100101",
 3779 => "00000010",
 3780 => "00111000",
 3781 => "00010101",
 3782 => "00101001",
 3783 => "00110100",
 3784 => "01010100",
 3785 => "11101100",
 3786 => "01000110",
 3787 => "10111001",
 3788 => "10000000",
 3789 => "00010001",
 3790 => "11011011",
 3791 => "10001000",
 3792 => "01011110",
 3793 => "01010101",
 3794 => "11100010",
 3795 => "10001110",
 3796 => "01001101",
 3797 => "10100010",
 3798 => "10100010",
 3799 => "00001101",
 3800 => "11111000",
 3801 => "00010100",
 3802 => "01011010",
 3803 => "11100101",
 3804 => "10000001",
 3805 => "10000011",
 3806 => "10010011",
 3807 => "01111011",
 3808 => "01000100",
 3809 => "11110101",
 3810 => "01100011",
 3811 => "00110010",
 3812 => "01101010",
 3813 => "11101111",
 3814 => "11111101",
 3815 => "00110001",
 3816 => "00000100",
 3817 => "11011100",
 3818 => "00100001",
 3819 => "01000100",
 3820 => "01010000",
 3821 => "11110010",
 3822 => "10100011",
 3823 => "10011110",
 3824 => "01010000",
 3825 => "10010111",
 3826 => "10111000",
 3827 => "10000110",
 3828 => "00101110",
 3829 => "11011110",
 3830 => "10000110",
 3831 => "10001001",
 3832 => "11110101",
 3833 => "01110001",
 3834 => "11110010",
 3835 => "01101100",
 3836 => "11001000",
 3837 => "10000001",
 3838 => "10010010",
 3839 => "10001110",
 3840 => "11100100",
 3841 => "00111101",
 3842 => "00010110",
 3843 => "00110001",
 3844 => "00010111",
 3845 => "00111001",
 3846 => "10011100",
 3847 => "00101010",
 3848 => "00110011",
 3849 => "10110111",
 3850 => "01010011",
 3851 => "10001110",
 3852 => "01110000",
 3853 => "00011101",
 3854 => "10001011",
 3855 => "01111011",
 3856 => "01010011",
 3857 => "00011000",
 3858 => "10101001",
 3859 => "01001010",
 3860 => "10111111",
 3861 => "01000011",
 3862 => "00011010",
 3863 => "00100000",
 3864 => "01111110",
 3865 => "00100101",
 3866 => "11011000",
 3867 => "11100011",
 3868 => "11111010",
 3869 => "00101100",
 3870 => "00001100",
 3871 => "01110000",
 3872 => "01100110",
 3873 => "10111000",
 3874 => "10110100",
 3875 => "10001110",
 3876 => "01011100",
 3877 => "11100011",
 3878 => "11111001",
 3879 => "10001000",
 3880 => "01110011",
 3881 => "01111111",
 3882 => "10110000",
 3883 => "10110011",
 3884 => "01001011",
 3885 => "10010011",
 3886 => "01110100",
 3887 => "01110000",
 3888 => "00011111",
 3889 => "10001001",
 3890 => "11101001",
 3891 => "00101010",
 3892 => "00000100",
 3893 => "10100111",
 3894 => "10101101",
 3895 => "01111111",
 3896 => "01101001",
 3897 => "10011001",
 3898 => "01000010",
 3899 => "00011101",
 3900 => "11011001",
 3901 => "11100010",
 3902 => "01110000",
 3903 => "11001110",
 3904 => "10101010",
 3905 => "11111111",
 3906 => "10011011",
 3907 => "01000101",
 3908 => "00001101",
 3909 => "11000100",
 3910 => "01111011",
 3911 => "01101000",
 3912 => "00101100",
 3913 => "01000000",
 3914 => "11101100",
 3915 => "11111001",
 3916 => "01001100",
 3917 => "11001111",
 3918 => "00111110",
 3919 => "00110100",
 3920 => "10101010",
 3921 => "11111100",
 3922 => "10011111",
 3923 => "01001100",
 3924 => "00010011",
 3925 => "00101101",
 3926 => "10110111",
 3927 => "10001011",
 3928 => "10110000",
 3929 => "00010011",
 3930 => "10000111",
 3931 => "01111001",
 3932 => "11010101",
 3933 => "10010111",
 3934 => "00001101",
 3935 => "11110001",
 3936 => "11011111",
 3937 => "01101001",
 3938 => "10110110",
 3939 => "00111100",
 3940 => "10101111",
 3941 => "10100001",
 3942 => "10001101",
 3943 => "01011100",
 3944 => "11101101",
 3945 => "01001001",
 3946 => "00111011",
 3947 => "01111011",
 3948 => "11010010",
 3949 => "00011110",
 3950 => "00010001",
 3951 => "01000000",
 3952 => "01001010",
 3953 => "10001000",
 3954 => "01110101",
 3955 => "10010100",
 3956 => "00001000",
 3957 => "11010000",
 3958 => "00010100",
 3959 => "10001101",
 3960 => "10101011",
 3961 => "10100100",
 3962 => "11101100",
 3963 => "10101111",
 3964 => "00101111",
 3965 => "11010111",
 3966 => "11111101",
 3967 => "10010101",
 3968 => "01000000",
 3969 => "01110011",
 3970 => "01111111",
 3971 => "01000001",
 3972 => "10110111",
 3973 => "10000110",
 3974 => "01010011",
 3975 => "11111100",
 3976 => "10000111",
 3977 => "00111110",
 3978 => "10010010",
 3979 => "01000000",
 3980 => "11101000",
 3981 => "11101001",
 3982 => "10000101",
 3983 => "11011011",
 3984 => "01001000",
 3985 => "10000010",
 3986 => "10110100",
 3987 => "11110010",
 3988 => "00011001",
 3989 => "10100001",
 3990 => "01010100",
 3991 => "11001101",
 3992 => "11010101",
 3993 => "11101111",
 3994 => "00100001",
 3995 => "00101001",
 3996 => "11100010",
 3997 => "11100010",
 3998 => "11011100",
 3999 => "10010011",
 4000 => "11010101",
 4001 => "01101101",
 4002 => "10011011",
 4003 => "01101100",
 4004 => "00010111",
 4005 => "10110110",
 4006 => "10110100",
 4007 => "00110111",
 4008 => "01010101",
 4009 => "11100100",
 4010 => "10101011",
 4011 => "11011001",
 4012 => "00101011",
 4013 => "10010000",
 4014 => "11110100",
 4015 => "11111000",
 4016 => "00000000",
 4017 => "01110000",
 4018 => "01111100",
 4019 => "11011001",
 4020 => "01000111",
 4021 => "00101010",
 4022 => "01101100",
 4023 => "10101101",
 4024 => "01100101",
 4025 => "11110011",
 4026 => "11010000",
 4027 => "01110100",
 4028 => "11110011",
 4029 => "11111001",
 4030 => "01001100",
 4031 => "00110011",
 4032 => "11110011",
 4033 => "01101000",
 4034 => "01011001",
 4035 => "01110111",
 4036 => "11110010",
 4037 => "01001111",
 4038 => "01111110",
 4039 => "01110111",
 4040 => "00011011",
 4041 => "11111010",
 4042 => "11001010",
 4043 => "00011010",
 4044 => "11001100",
 4045 => "11001111",
 4046 => "00111010",
 4047 => "00100110",
 4048 => "01011011",
 4049 => "10011010",
 4050 => "01110000",
 4051 => "10111011",
 4052 => "00111101",
 4053 => "11111111",
 4054 => "11000001",
 4055 => "10110101",
 4056 => "10010001",
 4057 => "11010111",
 4058 => "11001001",
 4059 => "10011001",
 4060 => "00100110",
 4061 => "10010111",
 4062 => "00110100",
 4063 => "01111100",
 4064 => "01011001",
 4065 => "00100011",
 4066 => "00100101",
 4067 => "10101111",
 4068 => "11101110",
 4069 => "00110100",
 4070 => "00000001",
 4071 => "10011010",
 4072 => "11100010",
 4073 => "10010100",
 4074 => "01011000",
 4075 => "01110111",
 4076 => "11100001",
 4077 => "11010111",
 4078 => "10110000",
 4079 => "00010011",
 4080 => "11101110",
 4081 => "10011100",
 4082 => "11101000",
 4083 => "01001110",
 4084 => "11011011",
 4085 => "01000100",
 4086 => "01111101",
 4087 => "11001110",
 4088 => "00000000",
 4089 => "00111111",
 4090 => "01011000",
 4091 => "00010000",
 4092 => "01100001",
 4093 => "00101110",
 4094 => "11010110",
 4095 => "01011000",
 4096 => "10110110",
 4097 => "00100110",
 4098 => "10100011",
 4099 => "11111111",
 4100 => "11011000",
 4101 => "10001100",
 4102 => "00010001",
 4103 => "01100100",
 4104 => "00000101",
 4105 => "00100010",
 4106 => "01101111",
 4107 => "01001101",
 4108 => "11111101",
 4109 => "01000011",
 4110 => "01001110",
 4111 => "00001010",
 4112 => "11001010",
 4113 => "10000111",
 4114 => "00010010",
 4115 => "01110001",
 4116 => "01100100",
 4117 => "01110000",
 4118 => "10101110",
 4119 => "11101101",
 4120 => "00011011",
 4121 => "10110011",
 4122 => "11110010",
 4123 => "00011000",
 4124 => "01110100",
 4125 => "01010000",
 4126 => "10101000",
 4127 => "11001101",
 4128 => "01001010",
 4129 => "10111001",
 4130 => "11110111",
 4131 => "11100111",
 4132 => "01001011",
 4133 => "01010001",
 4134 => "01010000",
 4135 => "11000101",
 4136 => "00111110",
 4137 => "00010110",
 4138 => "00000011",
 4139 => "10111010",
 4140 => "01100111",
 4141 => "00010101",
 4142 => "00101101",
 4143 => "11010010",
 4144 => "00001011",
 4145 => "10000100",
 4146 => "01001000",
 4147 => "11100001",
 4148 => "11111010",
 4149 => "01110001",
 4150 => "00011100",
 4151 => "11111100",
 4152 => "10101010",
 4153 => "01000000",
 4154 => "11101110",
 4155 => "01110111",
 4156 => "00010000",
 4157 => "00011100",
 4158 => "10000001",
 4159 => "10111011",
 4160 => "10000110",
 4161 => "01110101",
 4162 => "00111101",
 4163 => "00000010",
 4164 => "00101100",
 4165 => "00100111",
 4166 => "10011011",
 4167 => "10111011",
 4168 => "11011111",
 4169 => "01100101",
 4170 => "11110011",
 4171 => "11001011",
 4172 => "11001101",
 4173 => "01010101",
 4174 => "01100100",
 4175 => "00100011",
 4176 => "10101010",
 4177 => "11110100",
 4178 => "10110010",
 4179 => "11001100",
 4180 => "11110010",
 4181 => "11010010",
 4182 => "11111001",
 4183 => "10010011",
 4184 => "00110001",
 4185 => "11010000",
 4186 => "01101100",
 4187 => "10101010",
 4188 => "11110011",
 4189 => "11111011",
 4190 => "10111000",
 4191 => "11011110",
 4192 => "11111000",
 4193 => "00101101",
 4194 => "00100101",
 4195 => "10001000",
 4196 => "10110100",
 4197 => "01101010",
 4198 => "01011000",
 4199 => "11010000",
 4200 => "11110100",
 4201 => "01011001",
 4202 => "01100101",
 4203 => "11101111",
 4204 => "01110101",
 4205 => "00001111",
 4206 => "01001001",
 4207 => "00111111",
 4208 => "00111100",
 4209 => "10000100",
 4210 => "01111110",
 4211 => "11110100",
 4212 => "11101000",
 4213 => "10100110",
 4214 => "10001010",
 4215 => "01000000",
 4216 => "00000110",
 4217 => "00000111",
 4218 => "10000010",
 4219 => "01000010",
 4220 => "11111100",
 4221 => "00001101",
 4222 => "11001001",
 4223 => "00001110",
 4224 => "11111010",
 4225 => "11110001",
 4226 => "01010101",
 4227 => "00000110",
 4228 => "01101010",
 4229 => "00010100",
 4230 => "01101101",
 4231 => "01111001",
 4232 => "00111011",
 4233 => "11011100",
 4234 => "11010010",
 4235 => "10000100",
 4236 => "00011001",
 4237 => "01010011",
 4238 => "11110101",
 4239 => "11101000",
 4240 => "00000001",
 4241 => "01101010",
 4242 => "10101111",
 4243 => "01111011",
 4244 => "11110000",
 4245 => "10011111",
 4246 => "01000001",
 4247 => "01110000",
 4248 => "10011100",
 4249 => "11111001",
 4250 => "00011110",
 4251 => "00110000",
 4252 => "11001101",
 4253 => "01001111",
 4254 => "01100011",
 4255 => "01101001",
 4256 => "10101110",
 4257 => "10011000",
 4258 => "01010000",
 4259 => "00100101",
 4260 => "00010111",
 4261 => "10010010",
 4262 => "10101111",
 4263 => "10000000",
 4264 => "01010110",
 4265 => "11111010",
 4266 => "00010010",
 4267 => "01010011",
 4268 => "11110011",
 4269 => "11111010",
 4270 => "01010101",
 4271 => "00001001",
 4272 => "11001100",
 4273 => "01001100",
 4274 => "10010000",
 4275 => "11010100",
 4276 => "01011011",
 4277 => "00000110",
 4278 => "10100011",
 4279 => "00101001",
 4280 => "11011101",
 4281 => "11100011",
 4282 => "01000011",
 4283 => "00111101",
 4284 => "00000001",
 4285 => "10000000",
 4286 => "10001001",
 4287 => "10111010",
 4288 => "01001111",
 4289 => "11111101",
 4290 => "00001110",
 4291 => "01100110",
 4292 => "01111000",
 4293 => "10001000",
 4294 => "01011101",
 4295 => "10111001",
 4296 => "01110100",
 4297 => "10001010",
 4298 => "11101000",
 4299 => "00110100",
 4300 => "00101000",
 4301 => "01010101",
 4302 => "01000001",
 4303 => "10101100",
 4304 => "01000110",
 4305 => "00011000",
 4306 => "10101100",
 4307 => "00110100",
 4308 => "11101011",
 4309 => "10000101",
 4310 => "01011110",
 4311 => "00101011",
 4312 => "10011101",
 4313 => "10101111",
 4314 => "10111111",
 4315 => "01100101",
 4316 => "01000010",
 4317 => "10110001",
 4318 => "00010101",
 4319 => "00110010",
 4320 => "01111100",
 4321 => "01010010",
 4322 => "00110011",
 4323 => "01001111",
 4324 => "10101010",
 4325 => "00110110",
 4326 => "00110010",
 4327 => "11101011",
 4328 => "10001011",
 4329 => "01111101",
 4330 => "10100001",
 4331 => "11011100",
 4332 => "01101000",
 4333 => "01001000",
 4334 => "00111001",
 4335 => "01110010",
 4336 => "10111001",
 4337 => "01001010",
 4338 => "01101110",
 4339 => "00010001",
 4340 => "11011011",
 4341 => "10100001",
 4342 => "10001101",
 4343 => "11101111",
 4344 => "10110100",
 4345 => "10110110",
 4346 => "10010110",
 4347 => "11110101",
 4348 => "10011100",
 4349 => "10001100",
 4350 => "10101100",
 4351 => "10001111",
 4352 => "11110001",
 4353 => "11110000",
 4354 => "01011011",
 4355 => "00100100",
 4356 => "11101010",
 4357 => "10111011",
 4358 => "11010000",
 4359 => "01101011",
 4360 => "00100111",
 4361 => "11000001",
 4362 => "01101010",
 4363 => "10100011",
 4364 => "00100011",
 4365 => "00101010",
 4366 => "10101101",
 4367 => "00111001",
 4368 => "00001100",
 4369 => "00111010",
 4370 => "01111101",
 4371 => "10011010",
 4372 => "11111010",
 4373 => "00011100",
 4374 => "00011010",
 4375 => "11001011",
 4376 => "00011100",
 4377 => "10001110",
 4378 => "01001110",
 4379 => "00001000",
 4380 => "11111001",
 4381 => "11111100",
 4382 => "10011000",
 4383 => "00110100",
 4384 => "11100111",
 4385 => "10100101",
 4386 => "10110001",
 4387 => "00111110",
 4388 => "00011101",
 4389 => "10101101",
 4390 => "01011111",
 4391 => "00100011",
 4392 => "00101100",
 4393 => "11100100",
 4394 => "11101110",
 4395 => "10011111",
 4396 => "00010110",
 4397 => "11010100",
 4398 => "10111100",
 4399 => "00110110",
 4400 => "10011100",
 4401 => "01100101",
 4402 => "00010011",
 4403 => "11101000",
 4404 => "10000010",
 4405 => "01110111",
 4406 => "10000000",
 4407 => "01100110",
 4408 => "00001101",
 4409 => "10000101",
 4410 => "00000001",
 4411 => "00011111",
 4412 => "10010001",
 4413 => "10011100",
 4414 => "00101110",
 4415 => "10111111",
 4416 => "01110101",
 4417 => "01010011",
 4418 => "10101001",
 4419 => "10101101",
 4420 => "10011000",
 4421 => "10101011",
 4422 => "10100100",
 4423 => "01100110",
 4424 => "01101110",
 4425 => "01100000",
 4426 => "01110000",
 4427 => "10011011",
 4428 => "10101000",
 4429 => "11111010",
 4430 => "01110101",
 4431 => "00011100",
 4432 => "10100000",
 4433 => "00110110",
 4434 => "00101000",
 4435 => "11101101",
 4436 => "11010010",
 4437 => "01001110",
 4438 => "10001110",
 4439 => "11001000",
 4440 => "11111101",
 4441 => "11110110",
 4442 => "01101001",
 4443 => "11010010",
 4444 => "01100001",
 4445 => "01100100",
 4446 => "01000101",
 4447 => "01000110",
 4448 => "10000010",
 4449 => "00010101",
 4450 => "00100111",
 4451 => "01111110",
 4452 => "10111000",
 4453 => "01100100",
 4454 => "11001110",
 4455 => "01110010",
 4456 => "00010010",
 4457 => "01100000",
 4458 => "11011011",
 4459 => "10000000",
 4460 => "00011000",
 4461 => "11101001",
 4462 => "00110001",
 4463 => "00010100",
 4464 => "01000000",
 4465 => "10000110",
 4466 => "10101110",
 4467 => "01000000",
 4468 => "00111010",
 4469 => "11110101",
 4470 => "11100100",
 4471 => "10001011",
 4472 => "10100100",
 4473 => "00010011",
 4474 => "11100000",
 4475 => "11000101",
 4476 => "00111110",
 4477 => "00100001",
 4478 => "01001001",
 4479 => "10100110",
 4480 => "11001000",
 4481 => "01000010",
 4482 => "10010001",
 4483 => "11100000",
 4484 => "11101111",
 4485 => "11101001",
 4486 => "00111100",
 4487 => "01010011",
 4488 => "10111010",
 4489 => "11110001",
 4490 => "01111100",
 4491 => "00000010",
 4492 => "10101000",
 4493 => "10000101",
 4494 => "10110001",
 4495 => "01011001",
 4496 => "11010011",
 4497 => "00001110",
 4498 => "10001010",
 4499 => "11000100",
 4500 => "10001000",
 4501 => "00000100",
 4502 => "10001010",
 4503 => "01001011",
 4504 => "00110000",
 4505 => "10110011",
 4506 => "11110111",
 4507 => "11100111",
 4508 => "11111010",
 4509 => "10101000",
 4510 => "11010000",
 4511 => "10000011",
 4512 => "11101101",
 4513 => "01001100",
 4514 => "11000001",
 4515 => "10010010",
 4516 => "01111111",
 4517 => "01010110",
 4518 => "00001111",
 4519 => "00100101",
 4520 => "11111111",
 4521 => "11001110",
 4522 => "11111101",
 4523 => "11100101",
 4524 => "10010110",
 4525 => "11100100",
 4526 => "11001111",
 4527 => "11101100",
 4528 => "01010101",
 4529 => "10010100",
 4530 => "11011110",
 4531 => "00111101",
 4532 => "10010100",
 4533 => "00101101",
 4534 => "11011110",
 4535 => "00100111",
 4536 => "00000001",
 4537 => "01101010",
 4538 => "10000101",
 4539 => "10101000",
 4540 => "10001011",
 4541 => "10011111",
 4542 => "10010010",
 4543 => "01011010",
 4544 => "10001011",
 4545 => "01011011",
 4546 => "11111101",
 4547 => "10001010",
 4548 => "11011111",
 4549 => "00011000",
 4550 => "11000100",
 4551 => "10000101",
 4552 => "11001111",
 4553 => "10110010",
 4554 => "00100110",
 4555 => "00010111",
 4556 => "11001010",
 4557 => "11011011",
 4558 => "10110001",
 4559 => "01001100",
 4560 => "01110111",
 4561 => "10100110",
 4562 => "11101011",
 4563 => "01010001",
 4564 => "10110001",
 4565 => "00111100",
 4566 => "01111001",
 4567 => "11011111",
 4568 => "10001101",
 4569 => "00111010",
 4570 => "11010011",
 4571 => "00010110",
 4572 => "10000010",
 4573 => "10100101",
 4574 => "10101011",
 4575 => "10100110",
 4576 => "00100011",
 4577 => "10011010",
 4578 => "01101101",
 4579 => "01000001",
 4580 => "11101001",
 4581 => "01010111",
 4582 => "00101000",
 4583 => "11111001",
 4584 => "01101110",
 4585 => "10010100",
 4586 => "11111001",
 4587 => "00101100",
 4588 => "10000111",
 4589 => "00011110",
 4590 => "01110111",
 4591 => "01011110",
 4592 => "01001111",
 4593 => "10000000",
 4594 => "01101110",
 4595 => "01010011",
 4596 => "11111110",
 4597 => "10011011",
 4598 => "10111101",
 4599 => "11001110",
 4600 => "00011000",
 4601 => "10011100",
 4602 => "10110001",
 4603 => "01001001",
 4604 => "10111001",
 4605 => "01011000",
 4606 => "00000111",
 4607 => "11101010",
 4608 => "11101001",
 4609 => "11101010",
 4610 => "01010111",
 4611 => "10011001",
 4612 => "00111001",
 4613 => "01110000",
 4614 => "10101111",
 4615 => "01001110",
 4616 => "01000111",
 4617 => "11011101",
 4618 => "11011101",
 4619 => "00100110",
 4620 => "11011011",
 4621 => "10010100",
 4622 => "00100010",
 4623 => "01011000",
 4624 => "00011101",
 4625 => "11010101",
 4626 => "00000101",
 4627 => "10010000",
 4628 => "01110111",
 4629 => "10001001",
 4630 => "11000001",
 4631 => "10111010",
 4632 => "00110000",
 4633 => "11001001",
 4634 => "01000011",
 4635 => "11000110",
 4636 => "10101101",
 4637 => "11000110",
 4638 => "11100110",
 4639 => "01101101",
 4640 => "11101100",
 4641 => "01110011",
 4642 => "01100100",
 4643 => "01010011",
 4644 => "01011011",
 4645 => "10001111",
 4646 => "10101111",
 4647 => "00011011",
 4648 => "00011010",
 4649 => "00100101",
 4650 => "10001101",
 4651 => "01000010",
 4652 => "01011100",
 4653 => "11011010",
 4654 => "10110000",
 4655 => "11101100",
 4656 => "11000011",
 4657 => "11000100",
 4658 => "10100100",
 4659 => "11011111",
 4660 => "00001001",
 4661 => "00000100",
 4662 => "11111110",
 4663 => "00010101",
 4664 => "11010100",
 4665 => "01101001",
 4666 => "01111100",
 4667 => "11101000",
 4668 => "10010000",
 4669 => "01011010",
 4670 => "00101111",
 4671 => "11001001",
 4672 => "01110100",
 4673 => "10010001",
 4674 => "01001110",
 4675 => "10000101",
 4676 => "01000000",
 4677 => "11000110",
 4678 => "01110101",
 4679 => "11001100",
 4680 => "01011010",
 4681 => "11010001",
 4682 => "01010000",
 4683 => "11111000",
 4684 => "11010110",
 4685 => "00111010",
 4686 => "01011001",
 4687 => "11101001",
 4688 => "10100100",
 4689 => "01001011",
 4690 => "01100101",
 4691 => "11011011",
 4692 => "11110000",
 4693 => "01111110",
 4694 => "00000111",
 4695 => "01010101",
 4696 => "00101010",
 4697 => "11101010",
 4698 => "01100111",
 4699 => "01001101",
 4700 => "00101001",
 4701 => "00100101",
 4702 => "10100001",
 4703 => "01100001",
 4704 => "11011001",
 4705 => "10111100",
 4706 => "00011100",
 4707 => "11011110",
 4708 => "00100101",
 4709 => "01110110",
 4710 => "10110100",
 4711 => "01011110",
 4712 => "10010111",
 4713 => "10110010",
 4714 => "00001000",
 4715 => "01111101",
 4716 => "00101010",
 4717 => "01101111",
 4718 => "10000011",
 4719 => "11111101",
 4720 => "11110011",
 4721 => "01010001",
 4722 => "01011011",
 4723 => "01011000",
 4724 => "10011110",
 4725 => "11011111",
 4726 => "00000000",
 4727 => "00001011",
 4728 => "01101101",
 4729 => "00000000",
 4730 => "11101011",
 4731 => "00110010",
 4732 => "11000110",
 4733 => "00100101",
 4734 => "11000100",
 4735 => "11000101",
 4736 => "00000111",
 4737 => "10011101",
 4738 => "10001100",
 4739 => "00100010",
 4740 => "01001011",
 4741 => "00100011",
 4742 => "10001100",
 4743 => "10101010",
 4744 => "11010100",
 4745 => "01111101",
 4746 => "01000011",
 4747 => "10100011",
 4748 => "01011100",
 4749 => "01000101",
 4750 => "00100110",
 4751 => "01111110",
 4752 => "01010000",
 4753 => "11110011",
 4754 => "01001010",
 4755 => "00110101",
 4756 => "00000000",
 4757 => "01001010",
 4758 => "01011010",
 4759 => "11010010",
 4760 => "11111000",
 4761 => "10010110",
 4762 => "10111111",
 4763 => "10101010",
 4764 => "00100100",
 4765 => "11000100",
 4766 => "11000011",
 4767 => "00100101",
 4768 => "01101100",
 4769 => "10110011",
 4770 => "01010101",
 4771 => "11111111",
 4772 => "11000011",
 4773 => "11101111",
 4774 => "01110110",
 4775 => "00001110",
 4776 => "11101100",
 4777 => "00011111",
 4778 => "11110001",
 4779 => "01001010",
 4780 => "11011001",
 4781 => "00101101",
 4782 => "10100011",
 4783 => "00000011",
 4784 => "00111110",
 4785 => "00011101",
 4786 => "11111010",
 4787 => "10011010",
 4788 => "00000001",
 4789 => "00001101",
 4790 => "01011110",
 4791 => "01010110",
 4792 => "10111100",
 4793 => "01010011",
 4794 => "01100110",
 4795 => "10100011",
 4796 => "01010011",
 4797 => "10011100",
 4798 => "00001100",
 4799 => "00111011",
 4800 => "10100010",
 4801 => "10100110",
 4802 => "11011011",
 4803 => "11000001",
 4804 => "01001111",
 4805 => "01000010",
 4806 => "01100011",
 4807 => "01000110",
 4808 => "00100010",
 4809 => "11000110",
 4810 => "01001011",
 4811 => "11100011",
 4812 => "11101001",
 4813 => "00101000",
 4814 => "11110001",
 4815 => "01101001",
 4816 => "11110111",
 4817 => "10100110",
 4818 => "00001111",
 4819 => "00111011",
 4820 => "11100101",
 4821 => "00010011",
 4822 => "10111100",
 4823 => "00100011",
 4824 => "00001110",
 4825 => "01101010",
 4826 => "01110100",
 4827 => "10101000",
 4828 => "10001011",
 4829 => "00110110",
 4830 => "01000111",
 4831 => "10111011",
 4832 => "11011100",
 4833 => "01010110",
 4834 => "11100000",
 4835 => "00101010",
 4836 => "01100100",
 4837 => "00010011",
 4838 => "10010101",
 4839 => "00110011",
 4840 => "01000101",
 4841 => "10011000",
 4842 => "10011110",
 4843 => "11110001",
 4844 => "00000010",
 4845 => "01010011",
 4846 => "11011000",
 4847 => "01010001",
 4848 => "01111110",
 4849 => "00101001",
 4850 => "10001011",
 4851 => "10010011",
 4852 => "10011101",
 4853 => "00101111",
 4854 => "10001000",
 4855 => "00101110",
 4856 => "00000100",
 4857 => "00000010",
 4858 => "01010110",
 4859 => "10110100",
 4860 => "01100100",
 4861 => "00110100",
 4862 => "01100110",
 4863 => "01100100",
 4864 => "11100101",
 4865 => "11011100",
 4866 => "00011010",
 4867 => "00110101",
 4868 => "11101001",
 4869 => "10101011",
 4870 => "00111100",
 4871 => "10001001",
 4872 => "00101111",
 4873 => "00110001",
 4874 => "00100111",
 4875 => "11011110",
 4876 => "11001100",
 4877 => "11100101",
 4878 => "10001001",
 4879 => "10010100",
 4880 => "11010111",
 4881 => "00011111",
 4882 => "11111100",
 4883 => "11011001",
 4884 => "01110011",
 4885 => "10110010",
 4886 => "11100001",
 4887 => "11101101",
 4888 => "00110100",
 4889 => "01100110",
 4890 => "00100100",
 4891 => "11001111",
 4892 => "11111101",
 4893 => "01101101",
 4894 => "01010010",
 4895 => "10110011",
 4896 => "11001101",
 4897 => "10001111",
 4898 => "11011010",
 4899 => "01100110",
 4900 => "11000010",
 4901 => "11111010",
 4902 => "00001011",
 4903 => "10010110",
 4904 => "00100101",
 4905 => "00100010",
 4906 => "10110011",
 4907 => "10111110",
 4908 => "00111110",
 4909 => "00110011",
 4910 => "01001000",
 4911 => "00001000",
 4912 => "11110001",
 4913 => "00101001",
 4914 => "01011100",
 4915 => "00011100",
 4916 => "01101001",
 4917 => "11010000",
 4918 => "11000110",
 4919 => "00010010",
 4920 => "10001011",
 4921 => "10000000",
 4922 => "01011101",
 4923 => "00011011",
 4924 => "01101001",
 4925 => "11001010",
 4926 => "11011101",
 4927 => "00110010",
 4928 => "01010001",
 4929 => "01100100",
 4930 => "00001101",
 4931 => "11010110",
 4932 => "01011100",
 4933 => "10110101",
 4934 => "00000100",
 4935 => "00000110",
 4936 => "10100010",
 4937 => "11011101",
 4938 => "01011011",
 4939 => "10100111",
 4940 => "00001110",
 4941 => "01011110",
 4942 => "11100000",
 4943 => "00011001",
 4944 => "01010111",
 4945 => "10100011",
 4946 => "00110100",
 4947 => "10001000",
 4948 => "01000000",
 4949 => "10110011",
 4950 => "00000001",
 4951 => "00000101",
 4952 => "00101000",
 4953 => "11110100",
 4954 => "01010100",
 4955 => "01000011",
 4956 => "10110100",
 4957 => "01110100",
 4958 => "10010110",
 4959 => "01111110",
 4960 => "01111111",
 4961 => "10100000",
 4962 => "11001101",
 4963 => "11111001",
 4964 => "00100100",
 4965 => "10110110",
 4966 => "00110111",
 4967 => "01100101",
 4968 => "11101010",
 4969 => "00010010",
 4970 => "01001000",
 4971 => "11001010",
 4972 => "10100001",
 4973 => "00011010",
 4974 => "11101101",
 4975 => "00010111",
 4976 => "00000001",
 4977 => "11111000",
 4978 => "00011100",
 4979 => "11000110",
 4980 => "11100101",
 4981 => "01100111",
 4982 => "01110100",
 4983 => "10000111",
 4984 => "11111001",
 4985 => "00001101",
 4986 => "10011010",
 4987 => "00001001",
 4988 => "00110001",
 4989 => "10010000",
 4990 => "00101100",
 4991 => "11111011",
 4992 => "00000101",
 4993 => "01010010",
 4994 => "01010010",
 4995 => "10111110",
 4996 => "00000110",
 4997 => "00100011",
 4998 => "10000000",
 4999 => "00001010",
 5000 => "11011111",
 5001 => "11110100",
 5002 => "10010010",
 5003 => "01001100",
 5004 => "10001111",
 5005 => "01010001",
 5006 => "01101000",
 5007 => "00111011",
 5008 => "10111001",
 5009 => "11100011",
 5010 => "10001110",
 5011 => "00100100",
 5012 => "11010111",
 5013 => "11001001",
 5014 => "00111001",
 5015 => "10011001",
 5016 => "01111010",
 5017 => "10101011",
 5018 => "00001000",
 5019 => "11111001",
 5020 => "11111100",
 5021 => "11010010",
 5022 => "10010001",
 5023 => "01001000",
 5024 => "10001110",
 5025 => "00010011",
 5026 => "01011100",
 5027 => "10101100",
 5028 => "01000101",
 5029 => "01101011",
 5030 => "11110000",
 5031 => "10100000",
 5032 => "11000101",
 5033 => "10100001",
 5034 => "00111101",
 5035 => "00011001",
 5036 => "11010001",
 5037 => "11011011",
 5038 => "10111111",
 5039 => "00011001",
 5040 => "00100110",
 5041 => "00100100",
 5042 => "00100010",
 5043 => "00001010",
 5044 => "11111110",
 5045 => "00100110",
 5046 => "01100010",
 5047 => "11100111",
 5048 => "01110001",
 5049 => "01000011",
 5050 => "10010100",
 5051 => "01100000",
 5052 => "10001001",
 5053 => "00010000",
 5054 => "01011001",
 5055 => "01001101",
 5056 => "10001011",
 5057 => "10010000",
 5058 => "10111110",
 5059 => "01010000",
 5060 => "10001100",
 5061 => "01011101",
 5062 => "10110100",
 5063 => "01000101",
 5064 => "11010001",
 5065 => "01001101",
 5066 => "11101001",
 5067 => "00010000",
 5068 => "00011000",
 5069 => "11011010",
 5070 => "01010010",
 5071 => "01000000",
 5072 => "01011100",
 5073 => "00110110",
 5074 => "11011000",
 5075 => "10101011",
 5076 => "01110001",
 5077 => "11100010",
 5078 => "10010101",
 5079 => "00001011",
 5080 => "00001011",
 5081 => "01101010",
 5082 => "10110110",
 5083 => "11100000",
 5084 => "11100100",
 5085 => "10110001",
 5086 => "00101101",
 5087 => "10101100",
 5088 => "01011111",
 5089 => "10100110",
 5090 => "00101010",
 5091 => "11101100",
 5092 => "11001010",
 5093 => "11001001",
 5094 => "00000110",
 5095 => "01001111",
 5096 => "11000100",
 5097 => "11101001",
 5098 => "11000100",
 5099 => "10011100",
 5100 => "01100010",
 5101 => "11011011",
 5102 => "11111011",
 5103 => "00110010",
 5104 => "11100111",
 5105 => "11010011",
 5106 => "10110001",
 5107 => "00010010",
 5108 => "10101101",
 5109 => "00011000",
 5110 => "10011000",
 5111 => "11111110",
 5112 => "00110010",
 5113 => "00101011",
 5114 => "01001011",
 5115 => "01101011",
 5116 => "11111010",
 5117 => "11110000",
 5118 => "00010010",
 5119 => "01010101",
 5120 => "00001001",
 5121 => "10010110",
 5122 => "01101010",
 5123 => "11110110",
 5124 => "00000011",
 5125 => "00110111",
 5126 => "10010100",
 5127 => "11011101",
 5128 => "01111001",
 5129 => "01001110",
 5130 => "01010111",
 5131 => "10001011",
 5132 => "01100010",
 5133 => "01001111",
 5134 => "00111100",
 5135 => "11000111",
 5136 => "10010111",
 5137 => "10010111",
 5138 => "10010110",
 5139 => "10101100",
 5140 => "00010110",
 5141 => "00010100",
 5142 => "00011110",
 5143 => "01110001",
 5144 => "10011000",
 5145 => "11001110",
 5146 => "01100110",
 5147 => "00011111",
 5148 => "11111011",
 5149 => "11111101",
 5150 => "01111100",
 5151 => "10011001",
 5152 => "11110111",
 5153 => "01111010",
 5154 => "01010010",
 5155 => "00101100",
 5156 => "01100110",
 5157 => "11011000",
 5158 => "00110100",
 5159 => "00001010",
 5160 => "11111010",
 5161 => "10111100",
 5162 => "11110001",
 5163 => "01010000",
 5164 => "01101101",
 5165 => "01001000",
 5166 => "01011101",
 5167 => "01000100",
 5168 => "01000001",
 5169 => "10101100",
 5170 => "11000101",
 5171 => "01001111",
 5172 => "01101110",
 5173 => "00000011",
 5174 => "01110100",
 5175 => "00011110",
 5176 => "10011001",
 5177 => "11101011",
 5178 => "10110100",
 5179 => "00001000",
 5180 => "01010100",
 5181 => "11101010",
 5182 => "00111111",
 5183 => "10101100",
 5184 => "11110001",
 5185 => "11011110",
 5186 => "01001110",
 5187 => "00100010",
 5188 => "11101100",
 5189 => "01010100",
 5190 => "10011011",
 5191 => "11000111",
 5192 => "11111001",
 5193 => "10001010",
 5194 => "10001000",
 5195 => "10100011",
 5196 => "01011111",
 5197 => "10101000",
 5198 => "10101100",
 5199 => "11101111",
 5200 => "01110000",
 5201 => "01111001",
 5202 => "11110100",
 5203 => "01110111",
 5204 => "01011011",
 5205 => "11101011",
 5206 => "01011101",
 5207 => "01011011",
 5208 => "01011111",
 5209 => "00111011",
 5210 => "00101101",
 5211 => "11110000",
 5212 => "11010011",
 5213 => "10111101",
 5214 => "00001010",
 5215 => "11010110",
 5216 => "11101010",
 5217 => "11010100",
 5218 => "00110000",
 5219 => "11010100",
 5220 => "00100110",
 5221 => "00010001",
 5222 => "00101011",
 5223 => "01110001",
 5224 => "00100001",
 5225 => "11001110",
 5226 => "00101010",
 5227 => "01111101",
 5228 => "10101000",
 5229 => "00000101",
 5230 => "00101001",
 5231 => "00001010",
 5232 => "00111000",
 5233 => "10110110",
 5234 => "10100110",
 5235 => "11111110",
 5236 => "10011110",
 5237 => "11110110",
 5238 => "10011101",
 5239 => "11010100",
 5240 => "10100001",
 5241 => "10001110",
 5242 => "01111001",
 5243 => "10100001",
 5244 => "01101111",
 5245 => "11011101",
 5246 => "00001101",
 5247 => "10100011",
 5248 => "11001110",
 5249 => "10001111",
 5250 => "10111010",
 5251 => "01011101",
 5252 => "10100010",
 5253 => "10111111",
 5254 => "00000110",
 5255 => "01000111",
 5256 => "10110011",
 5257 => "00011010",
 5258 => "01000000",
 5259 => "11101110",
 5260 => "00011001",
 5261 => "01100101",
 5262 => "10101011",
 5263 => "01101111",
 5264 => "10110010",
 5265 => "01000011",
 5266 => "00101010",
 5267 => "01111110",
 5268 => "00100101",
 5269 => "11100010",
 5270 => "11101100",
 5271 => "10010100",
 5272 => "00111110",
 5273 => "10111001",
 5274 => "01111011",
 5275 => "01001011",
 5276 => "10010110",
 5277 => "11001100",
 5278 => "01101010",
 5279 => "11101001",
 5280 => "01001101",
 5281 => "10101001",
 5282 => "00111010",
 5283 => "10011100",
 5284 => "11111010",
 5285 => "10110001",
 5286 => "10000111",
 5287 => "00101010",
 5288 => "11110000",
 5289 => "11010111",
 5290 => "00000101",
 5291 => "10001001",
 5292 => "10110111",
 5293 => "01101010",
 5294 => "11000110",
 5295 => "01011011",
 5296 => "00111101",
 5297 => "00010010",
 5298 => "01000011",
 5299 => "11001100",
 5300 => "01000110",
 5301 => "11101001",
 5302 => "00001101",
 5303 => "00001000",
 5304 => "11000000",
 5305 => "10110010",
 5306 => "01000001",
 5307 => "10010011",
 5308 => "11100111",
 5309 => "00101010",
 5310 => "00011111",
 5311 => "11101101",
 5312 => "00001011",
 5313 => "10100101",
 5314 => "10001101",
 5315 => "10110001",
 5316 => "11011101",
 5317 => "01101101",
 5318 => "11000011",
 5319 => "00001111",
 5320 => "01101110",
 5321 => "10110001",
 5322 => "11100000",
 5323 => "10101010",
 5324 => "11111010",
 5325 => "00110110",
 5326 => "11000100",
 5327 => "01000000",
 5328 => "01101011",
 5329 => "00110010",
 5330 => "11000101",
 5331 => "10101100",
 5332 => "11100000",
 5333 => "11011101",
 5334 => "00101001",
 5335 => "01100001",
 5336 => "10110001",
 5337 => "00110010",
 5338 => "10001001",
 5339 => "10001000",
 5340 => "11000100",
 5341 => "11010110",
 5342 => "00001011",
 5343 => "10000101",
 5344 => "11011101",
 5345 => "10000100",
 5346 => "11001011",
 5347 => "10010011",
 5348 => "00011101",
 5349 => "00000111",
 5350 => "01111100",
 5351 => "00101101",
 5352 => "00001001",
 5353 => "11001111",
 5354 => "00101011",
 5355 => "11110101",
 5356 => "10010101",
 5357 => "00111110",
 5358 => "00111110",
 5359 => "00111100",
 5360 => "10111011",
 5361 => "01011001",
 5362 => "11100111",
 5363 => "00111011",
 5364 => "10110100",
 5365 => "00100000",
 5366 => "01100110",
 5367 => "00100110",
 5368 => "10001111",
 5369 => "10011111",
 5370 => "00011001",
 5371 => "01101001",
 5372 => "10001011",
 5373 => "00001100",
 5374 => "10010010",
 5375 => "00000110",
 5376 => "01001000",
 5377 => "11100101",
 5378 => "10000100",
 5379 => "00000101",
 5380 => "10011100",
 5381 => "11010001",
 5382 => "00011011",
 5383 => "11011100",
 5384 => "11010001",
 5385 => "11111001",
 5386 => "10111011",
 5387 => "01000111",
 5388 => "11011001",
 5389 => "01110100",
 5390 => "11011000",
 5391 => "01011100",
 5392 => "10110001",
 5393 => "10001100",
 5394 => "01100000",
 5395 => "01101111",
 5396 => "01111010",
 5397 => "01101011",
 5398 => "11000111",
 5399 => "00101101",
 5400 => "10011110",
 5401 => "10101100",
 5402 => "00010001",
 5403 => "00100011",
 5404 => "10100100",
 5405 => "00100011",
 5406 => "11100000",
 5407 => "10000010",
 5408 => "11100011",
 5409 => "01010101",
 5410 => "00111011",
 5411 => "11111010",
 5412 => "11010111",
 5413 => "10100010",
 5414 => "00111111",
 5415 => "00110011",
 5416 => "10001100",
 5417 => "01000101",
 5418 => "10101000",
 5419 => "00110010",
 5420 => "11010111",
 5421 => "10100011",
 5422 => "11101110",
 5423 => "01100110",
 5424 => "00100010",
 5425 => "10111100",
 5426 => "10010011",
 5427 => "11101111",
 5428 => "10111010",
 5429 => "00010011",
 5430 => "01110110",
 5431 => "10001010",
 5432 => "01000110",
 5433 => "00001111",
 5434 => "11000000",
 5435 => "00101111",
 5436 => "01111100",
 5437 => "00010010",
 5438 => "00011000",
 5439 => "11010000",
 5440 => "11100001",
 5441 => "00011111",
 5442 => "01010010",
 5443 => "10011101",
 5444 => "01110001",
 5445 => "01111011",
 5446 => "01100100",
 5447 => "10110011",
 5448 => "11010000",
 5449 => "00101100",
 5450 => "10001111",
 5451 => "11010010",
 5452 => "01001100",
 5453 => "10011011",
 5454 => "11111011",
 5455 => "11011100",
 5456 => "01100010",
 5457 => "00101100",
 5458 => "11110111",
 5459 => "00011011",
 5460 => "10011101",
 5461 => "01000100",
 5462 => "10101111",
 5463 => "10100111",
 5464 => "11001101",
 5465 => "10010111",
 5466 => "10111011",
 5467 => "01000011",
 5468 => "01101101",
 5469 => "01001100",
 5470 => "00010000",
 5471 => "00100110",
 5472 => "01101111",
 5473 => "11001111",
 5474 => "11101001",
 5475 => "01111101",
 5476 => "10111001",
 5477 => "01010010",
 5478 => "01101001",
 5479 => "01101011",
 5480 => "10000000",
 5481 => "00011110",
 5482 => "01111010",
 5483 => "11111100",
 5484 => "10000101",
 5485 => "00100101",
 5486 => "01111100",
 5487 => "00101010",
 5488 => "00001010",
 5489 => "01100011",
 5490 => "10011000",
 5491 => "00001011",
 5492 => "00001001",
 5493 => "00000001",
 5494 => "00011001",
 5495 => "01111111",
 5496 => "10001011",
 5497 => "00011110",
 5498 => "10110111",
 5499 => "11011111",
 5500 => "00110010",
 5501 => "10000011",
 5502 => "00001100",
 5503 => "10001011",
 5504 => "11100110",
 5505 => "10000000",
 5506 => "11110100",
 5507 => "01000100",
 5508 => "00100100",
 5509 => "10011000",
 5510 => "10101111",
 5511 => "01101000",
 5512 => "11111110",
 5513 => "01100111",
 5514 => "00011111",
 5515 => "01010100",
 5516 => "00000001",
 5517 => "11011110",
 5518 => "01011010",
 5519 => "00111000",
 5520 => "01100010",
 5521 => "01110010",
 5522 => "10011101",
 5523 => "00111110",
 5524 => "01011110",
 5525 => "10100101",
 5526 => "11111000",
 5527 => "01110010",
 5528 => "10100100",
 5529 => "01111000",
 5530 => "01100000",
 5531 => "10010001",
 5532 => "11111111",
 5533 => "10000110",
 5534 => "01000111",
 5535 => "11111001",
 5536 => "10100110",
 5537 => "01000100",
 5538 => "00101110",
 5539 => "01110001",
 5540 => "11110110",
 5541 => "10111111",
 5542 => "11001000",
 5543 => "00011110",
 5544 => "11011011",
 5545 => "10100001",
 5546 => "00111100",
 5547 => "00110011",
 5548 => "01000011",
 5549 => "01110010",
 5550 => "10100001",
 5551 => "11011011",
 5552 => "10110101",
 5553 => "00110100",
 5554 => "10010100",
 5555 => "11111001",
 5556 => "01101100",
 5557 => "00111010",
 5558 => "10010000",
 5559 => "10100101",
 5560 => "10000010",
 5561 => "10110110",
 5562 => "00010111",
 5563 => "01000010",
 5564 => "10101110",
 5565 => "01000110",
 5566 => "11011010",
 5567 => "00010111",
 5568 => "00100011",
 5569 => "00110110",
 5570 => "10100011",
 5571 => "10110110",
 5572 => "10100111",
 5573 => "11011000",
 5574 => "00101110",
 5575 => "01010001",
 5576 => "10010111",
 5577 => "11100000",
 5578 => "11110000",
 5579 => "11100101",
 5580 => "01011000",
 5581 => "00101100",
 5582 => "11111000",
 5583 => "10100101",
 5584 => "11101100",
 5585 => "01111001",
 5586 => "01000000",
 5587 => "10101010",
 5588 => "00011101",
 5589 => "10010100",
 5590 => "11100111",
 5591 => "01011101",
 5592 => "00011110",
 5593 => "01011110",
 5594 => "10011010",
 5595 => "10011100",
 5596 => "00101110",
 5597 => "00001011",
 5598 => "11101000",
 5599 => "00010000",
 5600 => "00100001",
 5601 => "00011010",
 5602 => "00010010",
 5603 => "00000101",
 5604 => "00111011",
 5605 => "11100100",
 5606 => "01011100",
 5607 => "10100000",
 5608 => "00010001",
 5609 => "11000011",
 5610 => "01001110",
 5611 => "11100100",
 5612 => "11100001",
 5613 => "01100001",
 5614 => "11110101",
 5615 => "01100110",
 5616 => "00101010",
 5617 => "00101000",
 5618 => "11110110",
 5619 => "10010001",
 5620 => "01111101",
 5621 => "00110100",
 5622 => "10100110",
 5623 => "10011100",
 5624 => "01010100",
 5625 => "00010000",
 5626 => "11000000",
 5627 => "00001100",
 5628 => "01001011",
 5629 => "01001110",
 5630 => "01001001",
 5631 => "10001111",
 5632 => "11011101",
 5633 => "10000010",
 5634 => "00001101",
 5635 => "01101110",
 5636 => "01010001",
 5637 => "11110100",
 5638 => "10001011",
 5639 => "01100000",
 5640 => "10010010",
 5641 => "00001011",
 5642 => "01101011",
 5643 => "11101010",
 5644 => "00010110",
 5645 => "01011100",
 5646 => "11011100",
 5647 => "10000101",
 5648 => "01010110",
 5649 => "11011000",
 5650 => "00011010",
 5651 => "10001111",
 5652 => "01001101",
 5653 => "11000001",
 5654 => "01111010",
 5655 => "01011011",
 5656 => "10100111",
 5657 => "11000011",
 5658 => "11011000",
 5659 => "00000100",
 5660 => "10100100",
 5661 => "11010000",
 5662 => "11011110",
 5663 => "01101010",
 5664 => "10001110",
 5665 => "10111001",
 5666 => "01111110",
 5667 => "01001101",
 5668 => "00001100",
 5669 => "01101001",
 5670 => "11110000",
 5671 => "10001010",
 5672 => "10000100",
 5673 => "11111100",
 5674 => "11110110",
 5675 => "11001100",
 5676 => "10010100",
 5677 => "11101100",
 5678 => "00101001",
 5679 => "11110000",
 5680 => "01110100",
 5681 => "10001001",
 5682 => "00110010",
 5683 => "10011011",
 5684 => "11001010",
 5685 => "10100101",
 5686 => "01011100",
 5687 => "10010110",
 5688 => "10100011",
 5689 => "01100111",
 5690 => "00111101",
 5691 => "01011110",
 5692 => "11011011",
 5693 => "10011101",
 5694 => "01011010",
 5695 => "10100000",
 5696 => "01011001",
 5697 => "01001001",
 5698 => "11010101",
 5699 => "00011101",
 5700 => "00100010",
 5701 => "11011000",
 5702 => "11001111",
 5703 => "01111011",
 5704 => "00000101",
 5705 => "10010010",
 5706 => "01100010",
 5707 => "11111001",
 5708 => "00001010",
 5709 => "10000111",
 5710 => "10000111",
 5711 => "10101100",
 5712 => "00000110",
 5713 => "00101001",
 5714 => "11010011",
 5715 => "11110111",
 5716 => "00100001",
 5717 => "10001010",
 5718 => "00111101",
 5719 => "00101000",
 5720 => "11110101",
 5721 => "01010100",
 5722 => "00000010",
 5723 => "01101001",
 5724 => "01000100",
 5725 => "00110111",
 5726 => "00101111",
 5727 => "10000111",
 5728 => "01000101",
 5729 => "11011100",
 5730 => "10101100",
 5731 => "00100101",
 5732 => "11100111",
 5733 => "01110101",
 5734 => "10010011",
 5735 => "10001100",
 5736 => "10011100",
 5737 => "11100000",
 5738 => "00110000",
 5739 => "00000110",
 5740 => "01001101",
 5741 => "01011000",
 5742 => "10010101",
 5743 => "00010111",
 5744 => "01111100",
 5745 => "11001001",
 5746 => "01000100",
 5747 => "10010011",
 5748 => "11100110",
 5749 => "00110100",
 5750 => "10011111",
 5751 => "01111111",
 5752 => "00101110",
 5753 => "01101110",
 5754 => "01100111",
 5755 => "01101101",
 5756 => "11110111",
 5757 => "11110111",
 5758 => "10101101",
 5759 => "01100110",
 5760 => "10010010",
 5761 => "11100010",
 5762 => "00100000",
 5763 => "01001011",
 5764 => "01110000",
 5765 => "01000110",
 5766 => "10001011",
 5767 => "11010001",
 5768 => "00000011",
 5769 => "10101001",
 5770 => "00000011",
 5771 => "10001111",
 5772 => "11100110",
 5773 => "01011000",
 5774 => "00010101",
 5775 => "01000011",
 5776 => "10110000",
 5777 => "00000101",
 5778 => "10011011",
 5779 => "11110011",
 5780 => "11100010",
 5781 => "01001110",
 5782 => "01000100",
 5783 => "10110010",
 5784 => "11000011",
 5785 => "00010110",
 5786 => "10110101",
 5787 => "01101101",
 5788 => "10001011",
 5789 => "10011001",
 5790 => "10100000",
 5791 => "10110001",
 5792 => "00010000",
 5793 => "11001100",
 5794 => "00010110",
 5795 => "01001011",
 5796 => "01011101",
 5797 => "11101011",
 5798 => "10011100",
 5799 => "11000100",
 5800 => "00111100",
 5801 => "10101110",
 5802 => "00000100",
 5803 => "01100101",
 5804 => "11000101",
 5805 => "01010000",
 5806 => "01001101",
 5807 => "00010101",
 5808 => "01011100",
 5809 => "11110000",
 5810 => "10011010",
 5811 => "11000010",
 5812 => "11101110",
 5813 => "00110000",
 5814 => "01011101",
 5815 => "01000000",
 5816 => "10011100",
 5817 => "01000101",
 5818 => "11101100",
 5819 => "01110110",
 5820 => "11111010",
 5821 => "10011110",
 5822 => "00110111",
 5823 => "11010000",
 5824 => "10011111",
 5825 => "01010111",
 5826 => "00000010",
 5827 => "11111011",
 5828 => "10011000",
 5829 => "11111011",
 5830 => "00000010",
 5831 => "11000011",
 5832 => "10010101",
 5833 => "00001010",
 5834 => "10001111",
 5835 => "00100100",
 5836 => "11011001",
 5837 => "01001000",
 5838 => "01100101",
 5839 => "10010000",
 5840 => "11111101",
 5841 => "10101001",
 5842 => "00001110",
 5843 => "10110010",
 5844 => "01111001",
 5845 => "11000001",
 5846 => "10001101",
 5847 => "10101110",
 5848 => "10101110",
 5849 => "11100000",
 5850 => "10000110",
 5851 => "00111101",
 5852 => "10100011",
 5853 => "01010111",
 5854 => "01100011",
 5855 => "00011011",
 5856 => "10100111",
 5857 => "11110000",
 5858 => "11101111",
 5859 => "01011110",
 5860 => "10000111",
 5861 => "10100011",
 5862 => "11001100",
 5863 => "10110101",
 5864 => "01000011",
 5865 => "00011111",
 5866 => "00011101",
 5867 => "10010001",
 5868 => "10111000",
 5869 => "10101010",
 5870 => "00001100",
 5871 => "01001000",
 5872 => "11000100",
 5873 => "01111000",
 5874 => "01101100",
 5875 => "00001101",
 5876 => "01110100",
 5877 => "01101111",
 5878 => "10001011",
 5879 => "10110011",
 5880 => "10111101",
 5881 => "11101011",
 5882 => "01010000",
 5883 => "11111110",
 5884 => "10011101",
 5885 => "01100110",
 5886 => "01011001",
 5887 => "10101001",
 5888 => "01100110",
 5889 => "10011011",
 5890 => "11001010",
 5891 => "11101000",
 5892 => "11010101",
 5893 => "10000110",
 5894 => "11010011",
 5895 => "01100110",
 5896 => "11001000",
 5897 => "11110101",
 5898 => "01101101",
 5899 => "01001001",
 5900 => "11101110",
 5901 => "00000011",
 5902 => "10011110",
 5903 => "10100111",
 5904 => "11011100",
 5905 => "10100101",
 5906 => "11100110",
 5907 => "10101000",
 5908 => "01010100",
 5909 => "10010110",
 5910 => "10110110",
 5911 => "01100110",
 5912 => "01111110",
 5913 => "01010011",
 5914 => "10000011",
 5915 => "10000110",
 5916 => "00110001",
 5917 => "01100010",
 5918 => "10010100",
 5919 => "11000110",
 5920 => "10100010",
 5921 => "11010111",
 5922 => "00111101",
 5923 => "10000001",
 5924 => "11000111",
 5925 => "10111000",
 5926 => "00001101",
 5927 => "00010001",
 5928 => "01101100",
 5929 => "11111110",
 5930 => "00110001",
 5931 => "10111010",
 5932 => "11000000",
 5933 => "00000100",
 5934 => "10101101",
 5935 => "11101000",
 5936 => "10111011",
 5937 => "00100101",
 5938 => "11001101",
 5939 => "00100010",
 5940 => "00001010",
 5941 => "10100110",
 5942 => "11101101",
 5943 => "00011011",
 5944 => "00111001",
 5945 => "11110011",
 5946 => "00011101",
 5947 => "10100110",
 5948 => "01100100",
 5949 => "11001010",
 5950 => "00000110",
 5951 => "11001110",
 5952 => "00110011",
 5953 => "00111101",
 5954 => "00111001",
 5955 => "01001000",
 5956 => "01000001",
 5957 => "00001100",
 5958 => "10101000",
 5959 => "11000111",
 5960 => "00000111",
 5961 => "01101101",
 5962 => "01100100",
 5963 => "01000100",
 5964 => "01011011",
 5965 => "10110110",
 5966 => "10011000",
 5967 => "01000100",
 5968 => "00011001",
 5969 => "10011111",
 5970 => "00101001",
 5971 => "11101100",
 5972 => "01100010",
 5973 => "00100100",
 5974 => "11101011",
 5975 => "11011010",
 5976 => "11001000",
 5977 => "11001100",
 5978 => "11100111",
 5979 => "10011010",
 5980 => "01001010",
 5981 => "10110111",
 5982 => "10101100",
 5983 => "11100110",
 5984 => "11010011",
 5985 => "00110101",
 5986 => "10011101",
 5987 => "00110101",
 5988 => "00000001",
 5989 => "11000000",
 5990 => "11100010",
 5991 => "01110110",
 5992 => "10110001",
 5993 => "10000011",
 5994 => "10111101",
 5995 => "11101100",
 5996 => "11100100",
 5997 => "00101011",
 5998 => "11010011",
 5999 => "00011110",
 6000 => "01010000",
 6001 => "00100011",
 6002 => "01000110",
 6003 => "00011101",
 6004 => "10100100",
 6005 => "11101101",
 6006 => "00110101",
 6007 => "10101001",
 6008 => "00001010",
 6009 => "10001000",
 6010 => "01011100",
 6011 => "00001100",
 6012 => "00000000",
 6013 => "01110110",
 6014 => "11011111",
 6015 => "00110110",
 6016 => "10111001",
 6017 => "11101011",
 6018 => "10111010",
 6019 => "10101110",
 6020 => "01001111",
 6021 => "00010111",
 6022 => "00101110",
 6023 => "11001001",
 6024 => "11000000",
 6025 => "00110100",
 6026 => "11011111",
 6027 => "01010011",
 6028 => "01110101",
 6029 => "10100100",
 6030 => "11100101",
 6031 => "10111000",
 6032 => "01000001",
 6033 => "01010000",
 6034 => "00010001",
 6035 => "00111011",
 6036 => "00111011",
 6037 => "00000010",
 6038 => "11100010",
 6039 => "01110000",
 6040 => "10100111",
 6041 => "00001101",
 6042 => "01011010",
 6043 => "01001000",
 6044 => "10101111",
 6045 => "10011101",
 6046 => "01011110",
 6047 => "00000100",
 6048 => "00010001",
 6049 => "10010010",
 6050 => "10101001",
 6051 => "00001100",
 6052 => "00000110",
 6053 => "00001001",
 6054 => "11111101",
 6055 => "10001100",
 6056 => "00101010",
 6057 => "00011111",
 6058 => "00001011",
 6059 => "11100100",
 6060 => "10110101",
 6061 => "00111000",
 6062 => "11110000",
 6063 => "11000000",
 6064 => "10111000",
 6065 => "10101110",
 6066 => "10000001",
 6067 => "01110100",
 6068 => "00001110",
 6069 => "10111101",
 6070 => "11111101",
 6071 => "10100011",
 6072 => "00011001",
 6073 => "01110001",
 6074 => "11100010",
 6075 => "10100100",
 6076 => "01100111",
 6077 => "00011100",
 6078 => "01101011",
 6079 => "10000111",
 6080 => "01110101",
 6081 => "10011010",
 6082 => "10010010",
 6083 => "11101000",
 6084 => "11110000",
 6085 => "00001110",
 6086 => "01110101",
 6087 => "11000001",
 6088 => "00111111",
 6089 => "11011010",
 6090 => "01101100",
 6091 => "01011100",
 6092 => "01011100",
 6093 => "10111000",
 6094 => "01100101",
 6095 => "00100101",
 6096 => "11000001",
 6097 => "00101001",
 6098 => "00110110",
 6099 => "11111111",
 6100 => "01101011",
 6101 => "10001111",
 6102 => "01101100",
 6103 => "11100100",
 6104 => "01010010",
 6105 => "00000001",
 6106 => "10010011",
 6107 => "11111110",
 6108 => "11111111",
 6109 => "11110110",
 6110 => "00011001",
 6111 => "11100110",
 6112 => "01011001",
 6113 => "00011011",
 6114 => "01001101",
 6115 => "00110001",
 6116 => "11110110",
 6117 => "00010111",
 6118 => "11001010",
 6119 => "10010000",
 6120 => "10111100",
 6121 => "01010000",
 6122 => "01001111",
 6123 => "00000010",
 6124 => "11101000",
 6125 => "01010001",
 6126 => "10100101",
 6127 => "11111110",
 6128 => "10000011",
 6129 => "00001000",
 6130 => "01000011",
 6131 => "11111010",
 6132 => "00101011",
 6133 => "00100111",
 6134 => "10000001",
 6135 => "00011111",
 6136 => "10011101",
 6137 => "00001111",
 6138 => "10010001",
 6139 => "10101101",
 6140 => "01000011",
 6141 => "10001111",
 6142 => "00100111",
 6143 => "00000011",
 6144 => "11110000",
 6145 => "01100111",
 6146 => "01011101",
 6147 => "01101011",
 6148 => "11011100",
 6149 => "11000110",
 6150 => "00111100",
 6151 => "11111010",
 6152 => "10100011",
 6153 => "11110001",
 6154 => "11011000",
 6155 => "11001001",
 6156 => "11001001",
 6157 => "11000011",
 6158 => "01011001",
 6159 => "01100101",
 6160 => "10001110",
 6161 => "10000111",
 6162 => "10001111",
 6163 => "00100111",
 6164 => "11110100",
 6165 => "11100000",
 6166 => "00010101",
 6167 => "11110001",
 6168 => "00000101",
 6169 => "10001111",
 6170 => "11100100",
 6171 => "01110010",
 6172 => "00000011",
 6173 => "10100100",
 6174 => "01100111",
 6175 => "00000111",
 6176 => "10100100",
 6177 => "10000010",
 6178 => "11010000",
 6179 => "11011110",
 6180 => "00001101",
 6181 => "00001110",
 6182 => "00111000",
 6183 => "01100010",
 6184 => "11011001",
 6185 => "00110100",
 6186 => "10100010",
 6187 => "01001011",
 6188 => "01101000",
 6189 => "11001101",
 6190 => "10111001",
 6191 => "11110001",
 6192 => "01101010",
 6193 => "11011001",
 6194 => "01000100",
 6195 => "11110010",
 6196 => "11100011",
 6197 => "11101110",
 6198 => "00011111",
 6199 => "10101001",
 6200 => "01100101",
 6201 => "11100100",
 6202 => "01110111",
 6203 => "00101100",
 6204 => "10011001",
 6205 => "10011101",
 6206 => "00101110",
 6207 => "01100000",
 6208 => "11111100",
 6209 => "10001111",
 6210 => "01001111",
 6211 => "01100011",
 6212 => "11110010",
 6213 => "01101011",
 6214 => "00010100",
 6215 => "11111100",
 6216 => "00001011",
 6217 => "01000100",
 6218 => "01010101",
 6219 => "00001010",
 6220 => "01111001",
 6221 => "00011110",
 6222 => "00111111",
 6223 => "10100110",
 6224 => "01111110",
 6225 => "00010001",
 6226 => "01100100",
 6227 => "00111010",
 6228 => "11101110",
 6229 => "01000100",
 6230 => "00100110",
 6231 => "10110111",
 6232 => "11010011",
 6233 => "10001001",
 6234 => "00011101",
 6235 => "11100100",
 6236 => "10111100",
 6237 => "00000110",
 6238 => "00101001",
 6239 => "10000101",
 6240 => "00001010",
 6241 => "10111100",
 6242 => "00101011",
 6243 => "00110011",
 6244 => "11101101",
 6245 => "10100110",
 6246 => "00111010",
 6247 => "10011000",
 6248 => "11001101",
 6249 => "11111001",
 6250 => "11111100",
 6251 => "00100110",
 6252 => "10010011",
 6253 => "10000000",
 6254 => "01011001",
 6255 => "11001110",
 6256 => "10011001",
 6257 => "01011011",
 6258 => "01111101",
 6259 => "11011000",
 6260 => "11110001",
 6261 => "10010111",
 6262 => "00000111",
 6263 => "01100000",
 6264 => "00000111",
 6265 => "01001010",
 6266 => "10011010",
 6267 => "10001111",
 6268 => "10101011",
 6269 => "01111101",
 6270 => "00010110",
 6271 => "01110111",
 6272 => "01001101",
 6273 => "00111001",
 6274 => "00000110",
 6275 => "01111110",
 6276 => "11000100",
 6277 => "10100011",
 6278 => "01110010",
 6279 => "00011000",
 6280 => "01010010",
 6281 => "00000100",
 6282 => "11001000",
 6283 => "11100011",
 6284 => "01000110",
 6285 => "10110101",
 6286 => "10000110",
 6287 => "01110110",
 6288 => "11010011",
 6289 => "01101000",
 6290 => "00100101",
 6291 => "11010011",
 6292 => "10101011",
 6293 => "11010000",
 6294 => "10101110",
 6295 => "11010101",
 6296 => "00011000",
 6297 => "01010011",
 6298 => "11010001",
 6299 => "00100010",
 6300 => "11101001",
 6301 => "01000110",
 6302 => "00110111",
 6303 => "01100111",
 6304 => "00010110",
 6305 => "00000001",
 6306 => "00000101",
 6307 => "00100001",
 6308 => "11100101",
 6309 => "11100100",
 6310 => "10100101",
 6311 => "01100101",
 6312 => "00111000",
 6313 => "11001110",
 6314 => "00001000",
 6315 => "01101011",
 6316 => "00010100",
 6317 => "11010101",
 6318 => "11111011",
 6319 => "00011000",
 6320 => "11010111",
 6321 => "01000100",
 6322 => "11110111",
 6323 => "11011101",
 6324 => "10000001",
 6325 => "11000101",
 6326 => "01001111",
 6327 => "01100001",
 6328 => "11010010",
 6329 => "01011001",
 6330 => "11001001",
 6331 => "11110010",
 6332 => "01111000",
 6333 => "11000001",
 6334 => "01111011",
 6335 => "00110101",
 6336 => "10011100",
 6337 => "10111100",
 6338 => "10100101",
 6339 => "01100100",
 6340 => "01001010",
 6341 => "01010101",
 6342 => "00110011",
 6343 => "10001010",
 6344 => "10100010",
 6345 => "01100111",
 6346 => "11001011",
 6347 => "00011001",
 6348 => "00011000",
 6349 => "10010001",
 6350 => "01101111",
 6351 => "00001011",
 6352 => "11010110",
 6353 => "11010000",
 6354 => "01011110",
 6355 => "00010110",
 6356 => "10100001",
 6357 => "11001110",
 6358 => "11001110",
 6359 => "11111100",
 6360 => "11110001",
 6361 => "00101111",
 6362 => "10001111",
 6363 => "00111011",
 6364 => "00000001",
 6365 => "11101111",
 6366 => "00101100",
 6367 => "10011001",
 6368 => "10011101",
 6369 => "10111110",
 6370 => "01010110",
 6371 => "01010110",
 6372 => "10010010",
 6373 => "01001100",
 6374 => "00000101",
 6375 => "01000111",
 6376 => "00110100",
 6377 => "11001001",
 6378 => "11111000",
 6379 => "01101100",
 6380 => "00111101",
 6381 => "11001101",
 6382 => "10110010",
 6383 => "01100111",
 6384 => "11011110",
 6385 => "00111101",
 6386 => "01000101",
 6387 => "11111000",
 6388 => "00100100",
 6389 => "00001101",
 6390 => "10000010",
 6391 => "10111100",
 6392 => "01000110",
 6393 => "01011111",
 6394 => "01100011",
 6395 => "11101000",
 6396 => "01001111",
 6397 => "11111001",
 6398 => "00000110",
 6399 => "01010100",
 6400 => "10010110",
 6401 => "01000100",
 6402 => "01010111",
 6403 => "01101010",
 6404 => "11000111",
 6405 => "00001101",
 6406 => "11010111",
 6407 => "00110111",
 6408 => "00001101",
 6409 => "10011100",
 6410 => "01110100",
 6411 => "10001111",
 6412 => "00000111",
 6413 => "10001011",
 6414 => "00011110",
 6415 => "01100000",
 6416 => "11011000",
 6417 => "10000010",
 6418 => "11010000",
 6419 => "00100000",
 6420 => "10010000",
 6421 => "10000110",
 6422 => "11111101",
 6423 => "11101100",
 6424 => "00110001",
 6425 => "01010110",
 6426 => "10101010",
 6427 => "01001010",
 6428 => "11010101",
 6429 => "00011000",
 6430 => "11101010",
 6431 => "10110110",
 6432 => "00110010",
 6433 => "00100110",
 6434 => "00010001",
 6435 => "11100100",
 6436 => "01100010",
 6437 => "00001000",
 6438 => "00100001",
 6439 => "10101010",
 6440 => "11010000",
 6441 => "00101011",
 6442 => "00111010",
 6443 => "11011110",
 6444 => "10110011",
 6445 => "10110101",
 6446 => "01101010",
 6447 => "00011100",
 6448 => "11110100",
 6449 => "11100100",
 6450 => "01010100",
 6451 => "00110110",
 6452 => "01111011",
 6453 => "01110000",
 6454 => "10111011",
 6455 => "10001010",
 6456 => "11111010",
 6457 => "11111001",
 6458 => "00101101",
 6459 => "10100100",
 6460 => "01111101",
 6461 => "10100111",
 6462 => "01111101",
 6463 => "00100011",
 6464 => "10100001",
 6465 => "11001011",
 6466 => "00101000",
 6467 => "10001010",
 6468 => "10000000",
 6469 => "01010110",
 6470 => "01100001",
 6471 => "01101000",
 6472 => "01000101",
 6473 => "10100010",
 6474 => "01000001",
 6475 => "01101010",
 6476 => "11110100",
 6477 => "11110110",
 6478 => "01110100",
 6479 => "00011001",
 6480 => "01001010",
 6481 => "11010100",
 6482 => "11100110",
 6483 => "10000000",
 6484 => "10000111",
 6485 => "11111101",
 6486 => "01011011",
 6487 => "00011111",
 6488 => "00000111",
 6489 => "00111000",
 6490 => "00110110",
 6491 => "01100011",
 6492 => "10111111",
 6493 => "00110011",
 6494 => "10001010",
 6495 => "10100110",
 6496 => "01000101",
 6497 => "10101001",
 6498 => "10101110",
 6499 => "11010101",
 6500 => "01101101",
 6501 => "01100100",
 6502 => "11001110",
 6503 => "01011101",
 6504 => "11011111", others => (others =>'0'));
component project_reti_logiche is 
    port (
            i_clk         : in  std_logic;
            i_start       : in  std_logic;
            i_rst         : in  std_logic;
            i_data       : in  std_logic_vector(7 downto 0); --1 byte
            o_address     : out std_logic_vector(15 downto 0); --16 bit addr: max size is 255*255 + 3 more for max x and y and thresh.
            o_done            : out std_logic;
            o_en         : out std_logic;
            o_we       : out std_logic;
            o_data            : out std_logic_vector (7 downto 0)
          );
end component project_reti_logiche;
begin 
	UUT: project_reti_logiche
	port map (
		  i_clk      	=> tb_clk,	
          i_start       => tb_start,
          i_rst      	=> tb_rst,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address, 
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
		  o_we 	=> mem_we,
          o_data    => mem_i_data
);p_CLK_GEN : process is
  begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
  end process p_CLK_GEN; 
 MEM : process(tb_clk)
   begin
    if tb_clk'event and tb_clk = '1' then
     if enable_wire = '1' then
      if mem_we = '1' then
       RAM(conv_integer(mem_address))              <= mem_i_data;
       mem_o_data                      <= mem_i_data;
      else
       mem_o_data <= RAM(conv_integer(mem_address));
      end if;
     end if;
    end if;
   end process;
test : process is
begin 
wait for 100 ns;
wait for c_CLOCK_PERIOD;
tb_rst <= '1';
wait for c_CLOCK_PERIOD;
tb_rst <= '0';
wait for c_CLOCK_PERIOD;
tb_start <= '1';
wait for c_CLOCK_PERIOD; 
tb_start <= '0';
wait until tb_done = '1';
wait until tb_done = '0';
wait until rising_edge(tb_clk);

 
assert RAM(1) = "00011001" report "FAIL high bits" severity failure;
assert RAM(0) = "01100100" report "FAIL low bits" severity failure;
assert false report "Simulation Ended!, test passed" severity failure;
end process test;
 end projecttb;