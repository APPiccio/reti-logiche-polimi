library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity project_tb is
end project_tb;
architecture projecttb of project_tb is
constant c_CLOCK_PERIOD		: time := 15 ns;
signal   tb_done		: std_logic;
signal   mem_address		: std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst		    : std_logic := '0';
signal   tb_start		: std_logic := '0';
signal   tb_clk		    : std_logic := '0';
signal   mem_o_data,mem_i_data		: std_logic_vector (7 downto 0);
signal   enable_wire  		: std_logic;
signal   mem_we		: std_logic;
type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
signal RAM: ram_type := (2 => "01000101", 3 => "10011110", 4 => "00011011",
 5 => "01010001",
 6 => "01110100",
 7 => "10011000",
 8 => "11110010",
 9 => "00011000",
 10 => "10101011",
 11 => "11111000",
 12 => "00100100",
 13 => "10101101",
 14 => "10001011",
 15 => "11100110",
 16 => "11001100",
 17 => "11111000",
 18 => "01110001",
 19 => "11010110",
 20 => "11100101",
 21 => "01111110",
 22 => "11101001",
 23 => "00100011",
 24 => "01001110",
 25 => "10011100",
 26 => "10111011",
 27 => "01010001",
 28 => "01011101",
 29 => "00100111",
 30 => "01110000",
 31 => "00101100",
 32 => "01110001",
 33 => "00111110",
 34 => "11101010",
 35 => "00000001",
 36 => "01010100",
 37 => "11001001",
 38 => "11011011",
 39 => "11100000",
 40 => "10001111",
 41 => "00110100",
 42 => "11100111",
 43 => "11010010",
 44 => "10010000",
 45 => "01010110",
 46 => "10010100",
 47 => "00000101",
 48 => "00100111",
 49 => "00010010",
 50 => "00000100",
 51 => "10000101",
 52 => "01010011",
 53 => "11111110",
 54 => "10010111",
 55 => "10101000",
 56 => "10000001",
 57 => "01010010",
 58 => "11110010",
 59 => "11101001",
 60 => "00100001",
 61 => "01011100",
 62 => "01010100",
 63 => "11111001",
 64 => "00100111",
 65 => "01010000",
 66 => "00101100",
 67 => "11100101",
 68 => "00000011",
 69 => "00001110",
 70 => "11100110",
 71 => "01110010",
 72 => "01001000",
 73 => "10001010",
 74 => "11110110",
 75 => "01001110",
 76 => "10000000",
 77 => "11011110",
 78 => "11010100",
 79 => "11101111",
 80 => "10000101",
 81 => "10100100",
 82 => "10010101",
 83 => "10001110",
 84 => "11000011",
 85 => "00111110",
 86 => "00011101",
 87 => "00111011",
 88 => "01101111",
 89 => "10011101",
 90 => "10100111",
 91 => "01010110",
 92 => "00101110",
 93 => "01001111",
 94 => "00101010",
 95 => "00000100",
 96 => "01110010",
 97 => "01001000",
 98 => "11010110",
 99 => "01100110",
 100 => "01000010",
 101 => "00111001",
 102 => "01110000",
 103 => "11011001",
 104 => "01110101",
 105 => "10101101",
 106 => "11110111",
 107 => "00010101",
 108 => "01110000",
 109 => "11001111",
 110 => "10110010",
 111 => "10011111",
 112 => "01101110",
 113 => "10110100",
 114 => "11010001",
 115 => "11101101",
 116 => "11010101",
 117 => "11011100",
 118 => "00010010",
 119 => "00100000",
 120 => "01110000",
 121 => "01001111",
 122 => "11011011",
 123 => "00100011",
 124 => "11010011",
 125 => "11100011",
 126 => "11010111",
 127 => "00010000",
 128 => "10011001",
 129 => "00011010",
 130 => "10001000",
 131 => "01111101",
 132 => "10101010",
 133 => "10000110",
 134 => "10110100",
 135 => "10010101",
 136 => "10010011",
 137 => "10000001",
 138 => "10000001",
 139 => "10001100",
 140 => "11001100",
 141 => "10011100",
 142 => "00000001",
 143 => "11101110",
 144 => "00111001",
 145 => "11010000",
 146 => "01001101",
 147 => "11100011",
 148 => "01100001",
 149 => "11100001",
 150 => "10000010",
 151 => "01100111",
 152 => "11100011",
 153 => "11001101",
 154 => "10011010",
 155 => "11111010",
 156 => "01111111",
 157 => "11100011",
 158 => "00001000",
 159 => "11000111",
 160 => "00100100",
 161 => "01111100",
 162 => "10011010",
 163 => "11001011",
 164 => "00100011",
 165 => "10111000",
 166 => "10110010",
 167 => "00101011",
 168 => "00000011",
 169 => "00010011",
 170 => "11000111",
 171 => "10010001",
 172 => "11100110",
 173 => "01001001",
 174 => "11100100",
 175 => "01101110",
 176 => "10000100",
 177 => "00000001",
 178 => "01110011",
 179 => "11100111",
 180 => "00111000",
 181 => "10010101",
 182 => "10100100",
 183 => "11101011",
 184 => "01011110",
 185 => "10011100",
 186 => "10011110",
 187 => "10111001",
 188 => "10011001",
 189 => "11001110",
 190 => "00000001",
 191 => "00110101",
 192 => "11011110",
 193 => "10100011",
 194 => "00011011",
 195 => "00111011",
 196 => "11100100",
 197 => "10101011",
 198 => "11001110",
 199 => "01000101",
 200 => "01011110",
 201 => "11111011",
 202 => "11010010",
 203 => "01110010",
 204 => "01000101",
 205 => "10011000",
 206 => "11000001",
 207 => "11111000",
 208 => "11100011",
 209 => "00101011",
 210 => "10100111",
 211 => "00111100",
 212 => "10100000",
 213 => "01101000",
 214 => "11000011",
 215 => "10001010",
 216 => "11110000",
 217 => "01101011",
 218 => "00111101",
 219 => "10111000",
 220 => "10000101",
 221 => "00101110",
 222 => "01101101",
 223 => "01011001",
 224 => "11001010",
 225 => "00111000",
 226 => "00001011",
 227 => "00101111",
 228 => "10110010",
 229 => "11000111",
 230 => "01010010",
 231 => "00010011",
 232 => "00000101",
 233 => "01111110",
 234 => "10010100",
 235 => "01100101",
 236 => "00000001",
 237 => "10000000",
 238 => "00110100",
 239 => "00110001",
 240 => "01011100",
 241 => "01100111",
 242 => "10011100",
 243 => "10110100",
 244 => "10101111",
 245 => "10000100",
 246 => "01111011",
 247 => "11111110",
 248 => "10010011",
 249 => "00010110",
 250 => "00011101",
 251 => "10100111",
 252 => "01101110",
 253 => "10101111",
 254 => "01001100",
 255 => "01110101",
 256 => "00010100",
 257 => "10010011",
 258 => "10011100",
 259 => "01010110",
 260 => "11010001",
 261 => "10010101",
 262 => "10111110",
 263 => "00001100",
 264 => "10101100",
 265 => "00001011",
 266 => "01011110",
 267 => "10110010",
 268 => "10110101",
 269 => "10100010",
 270 => "10101100",
 271 => "11101000",
 272 => "00110110",
 273 => "11110110",
 274 => "01101000",
 275 => "11010011",
 276 => "10010111",
 277 => "10101111",
 278 => "00011001",
 279 => "00101111",
 280 => "10000000",
 281 => "11000111",
 282 => "00110010",
 283 => "00000110",
 284 => "00110110",
 285 => "10000011",
 286 => "11111100",
 287 => "01111100",
 288 => "01000000",
 289 => "00110101",
 290 => "10011100",
 291 => "01111100",
 292 => "10001000",
 293 => "10100010",
 294 => "00001100",
 295 => "00011110",
 296 => "11100001",
 297 => "01111111",
 298 => "11100111",
 299 => "11100110",
 300 => "00000101",
 301 => "10000010",
 302 => "00101111",
 303 => "10110110",
 304 => "00001010",
 305 => "10000000",
 306 => "11011111",
 307 => "11110101",
 308 => "00101101",
 309 => "11101010",
 310 => "11110001",
 311 => "01000000",
 312 => "10010011",
 313 => "11110101",
 314 => "11110111",
 315 => "01101110",
 316 => "00011011",
 317 => "10011101",
 318 => "01011100",
 319 => "10100100",
 320 => "01001011",
 321 => "10100111",
 322 => "10000101",
 323 => "10111100",
 324 => "11001100",
 325 => "01100010",
 326 => "00101100",
 327 => "00101011",
 328 => "10011011",
 329 => "00010000",
 330 => "00100111",
 331 => "00111001",
 332 => "01011101",
 333 => "01010100",
 334 => "01101111",
 335 => "10001101",
 336 => "10010110",
 337 => "11001111",
 338 => "00000111",
 339 => "01111100",
 340 => "11101011",
 341 => "00101001",
 342 => "10100010",
 343 => "10100100",
 344 => "01010010",
 345 => "01111100",
 346 => "10110111",
 347 => "10001101",
 348 => "01001100",
 349 => "00010001",
 350 => "10010100",
 351 => "00010010",
 352 => "10011001",
 353 => "01101000",
 354 => "01001000",
 355 => "10011111",
 356 => "11111001",
 357 => "11000011",
 358 => "11100100",
 359 => "11111001",
 360 => "01101000",
 361 => "10110010",
 362 => "11001010",
 363 => "11101101",
 364 => "11011001",
 365 => "01100100",
 366 => "01010101",
 367 => "00111100",
 368 => "00101111",
 369 => "11111000",
 370 => "00111011",
 371 => "00001100",
 372 => "10101000",
 373 => "11101110",
 374 => "10111011",
 375 => "11000101",
 376 => "00010000",
 377 => "11010011",
 378 => "10101100",
 379 => "01000111",
 380 => "01101100",
 381 => "10011011",
 382 => "01100001",
 383 => "10101101",
 384 => "10110111",
 385 => "00010100",
 386 => "01011101",
 387 => "00100010",
 388 => "11011101",
 389 => "10011101",
 390 => "01001110",
 391 => "00101001",
 392 => "00010001",
 393 => "10111100",
 394 => "01110101",
 395 => "10010101",
 396 => "00001100",
 397 => "10010011",
 398 => "11111000",
 399 => "01110101",
 400 => "10010100",
 401 => "01011010",
 402 => "01110100",
 403 => "00100000",
 404 => "10110011",
 405 => "01101100",
 406 => "01110111",
 407 => "11110110",
 408 => "10100100",
 409 => "01000000",
 410 => "11010110",
 411 => "00001101",
 412 => "10000100",
 413 => "01011010",
 414 => "00000010",
 415 => "01010011",
 416 => "10111101",
 417 => "01101001",
 418 => "00111010",
 419 => "00011100",
 420 => "00000001",
 421 => "11101011",
 422 => "00101001",
 423 => "11001101",
 424 => "00101111",
 425 => "01001000",
 426 => "11010111",
 427 => "11110011",
 428 => "11111111",
 429 => "10011101",
 430 => "00010011",
 431 => "00011111",
 432 => "01000011",
 433 => "10101000",
 434 => "10111110",
 435 => "11001011",
 436 => "00001010",
 437 => "01100000",
 438 => "01011100",
 439 => "10101101",
 440 => "01100101",
 441 => "00100001",
 442 => "00100010",
 443 => "00001111",
 444 => "01000011",
 445 => "10001000",
 446 => "11011011",
 447 => "01010111",
 448 => "11000001",
 449 => "01000000",
 450 => "00010001",
 451 => "11010010",
 452 => "11010001",
 453 => "10010101",
 454 => "11000110",
 455 => "01011110",
 456 => "01001011",
 457 => "00010010",
 458 => "11001101",
 459 => "00110101",
 460 => "01101001",
 461 => "00011000",
 462 => "00101111",
 463 => "10000110",
 464 => "01000111",
 465 => "00010110",
 466 => "00001010",
 467 => "01001001",
 468 => "00110100",
 469 => "00111000",
 470 => "11011100",
 471 => "00110111",
 472 => "00111100",
 473 => "11010111",
 474 => "00000100",
 475 => "10110101",
 476 => "01011110",
 477 => "10011010",
 478 => "11110000",
 479 => "11010111",
 480 => "00011110",
 481 => "01000011",
 482 => "00101000",
 483 => "00101000",
 484 => "00011011",
 485 => "00110100",
 486 => "11010111",
 487 => "01000000",
 488 => "00100000",
 489 => "01001111",
 490 => "11011101",
 491 => "10100010",
 492 => "10011011",
 493 => "00100011",
 494 => "00111001",
 495 => "10011001",
 496 => "10001011",
 497 => "00100110",
 498 => "10010100",
 499 => "01100111",
 500 => "00100010",
 501 => "00101000",
 502 => "10101101",
 503 => "11001011",
 504 => "00000000",
 505 => "01110000",
 506 => "11011000",
 507 => "00001111",
 508 => "00010000",
 509 => "10101000",
 510 => "10010101",
 511 => "10010110",
 512 => "11001010",
 513 => "11110101",
 514 => "11101100",
 515 => "01111111",
 516 => "01111011",
 517 => "00100010",
 518 => "00101011",
 519 => "11001111",
 520 => "00100110",
 521 => "10010011",
 522 => "01100110",
 523 => "11100111",
 524 => "01000100",
 525 => "11100101",
 526 => "10110111",
 527 => "11110001",
 528 => "11100010",
 529 => "01100110",
 530 => "00111110",
 531 => "01111011",
 532 => "01000011",
 533 => "11101101",
 534 => "10101010",
 535 => "00010110",
 536 => "10010110",
 537 => "11111111",
 538 => "11001011",
 539 => "01111111",
 540 => "01011110",
 541 => "01001011",
 542 => "10111101",
 543 => "00001100",
 544 => "00101111",
 545 => "01111001",
 546 => "10001011",
 547 => "00101001",
 548 => "10000011",
 549 => "01000010",
 550 => "01111001",
 551 => "10110100",
 552 => "10111000",
 553 => "00001001",
 554 => "00110101",
 555 => "00111100",
 556 => "01111100",
 557 => "11001101",
 558 => "00111011",
 559 => "01110100",
 560 => "11000000",
 561 => "01101010",
 562 => "11000001",
 563 => "10110011",
 564 => "00110100",
 565 => "01101000",
 566 => "01000101",
 567 => "01100000",
 568 => "00111011",
 569 => "01110001",
 570 => "11100000",
 571 => "00111001",
 572 => "01110000",
 573 => "10000010",
 574 => "00000001",
 575 => "00000001",
 576 => "10010011",
 577 => "10111100",
 578 => "10110101",
 579 => "11001001",
 580 => "10000010",
 581 => "00010111",
 582 => "10010100",
 583 => "11010001",
 584 => "11100000",
 585 => "11011110",
 586 => "01110101",
 587 => "10100000",
 588 => "10010100",
 589 => "10101001",
 590 => "00110011",
 591 => "11000001",
 592 => "01000010",
 593 => "01110111",
 594 => "10011010",
 595 => "01111111",
 596 => "00001110",
 597 => "10111010",
 598 => "11111000",
 599 => "11001010",
 600 => "00100101",
 601 => "10100111",
 602 => "10001011",
 603 => "11111110",
 604 => "10010101",
 605 => "00000110",
 606 => "11001110",
 607 => "00000100",
 608 => "10110100",
 609 => "10010111",
 610 => "10100011",
 611 => "01111101",
 612 => "11000101",
 613 => "00001010",
 614 => "11100111",
 615 => "01000011",
 616 => "01000010",
 617 => "01100100",
 618 => "00111010",
 619 => "01111100",
 620 => "00110111",
 621 => "01011110",
 622 => "11000110",
 623 => "00101111",
 624 => "11111110",
 625 => "11010110",
 626 => "10100001",
 627 => "00001100",
 628 => "11000110",
 629 => "01001000",
 630 => "11010111",
 631 => "00111101",
 632 => "01110100",
 633 => "10011110",
 634 => "10101010",
 635 => "00110010",
 636 => "10000110",
 637 => "00011100",
 638 => "01001001",
 639 => "00001100",
 640 => "00101100",
 641 => "10101000",
 642 => "10110001",
 643 => "10001001",
 644 => "10111100",
 645 => "11100000",
 646 => "00000110",
 647 => "10001000",
 648 => "00111011",
 649 => "01010111",
 650 => "00111001",
 651 => "11001001",
 652 => "00001000",
 653 => "00100001",
 654 => "00001101",
 655 => "00111011",
 656 => "10100101",
 657 => "10010100",
 658 => "11111010",
 659 => "00011000",
 660 => "01100110",
 661 => "10011111",
 662 => "11010101",
 663 => "10001001",
 664 => "00101001",
 665 => "00100111",
 666 => "11111100",
 667 => "11011000",
 668 => "00111101",
 669 => "00111101",
 670 => "00001101",
 671 => "11101000",
 672 => "01001100",
 673 => "00010111",
 674 => "11110100",
 675 => "11011110",
 676 => "10000011",
 677 => "10111000",
 678 => "10110011",
 679 => "01001000",
 680 => "01011101",
 681 => "01010101",
 682 => "10100101",
 683 => "00001110",
 684 => "11000101",
 685 => "00001000",
 686 => "01001001",
 687 => "10111101",
 688 => "11001101",
 689 => "10001000",
 690 => "11101101",
 691 => "01100101",
 692 => "00100111",
 693 => "01001111",
 694 => "01110000",
 695 => "01001011",
 696 => "01011111",
 697 => "10010110",
 698 => "10010011",
 699 => "11011100",
 700 => "10100101",
 701 => "11110010",
 702 => "10010111",
 703 => "10011111",
 704 => "10111001",
 705 => "01101010",
 706 => "10111010",
 707 => "01111001",
 708 => "00101010",
 709 => "01101011",
 710 => "11000100",
 711 => "00101110",
 712 => "01001100",
 713 => "01100000",
 714 => "10100110",
 715 => "01111011",
 716 => "00100001",
 717 => "11011011",
 718 => "11001011",
 719 => "00111101",
 720 => "00111001",
 721 => "11000110",
 722 => "10001011",
 723 => "00011010",
 724 => "00010010",
 725 => "11101100",
 726 => "01101000",
 727 => "10001101",
 728 => "00011000",
 729 => "01110010",
 730 => "00011010",
 731 => "11011100",
 732 => "10000001",
 733 => "10001111",
 734 => "00000101",
 735 => "01000000",
 736 => "11011000",
 737 => "00101111",
 738 => "10000100",
 739 => "11000110",
 740 => "10100100",
 741 => "10101011",
 742 => "10011100",
 743 => "11110111",
 744 => "01001001",
 745 => "11010101",
 746 => "01101110",
 747 => "01101001",
 748 => "00000101",
 749 => "11111111",
 750 => "01001101",
 751 => "00101010",
 752 => "10011110",
 753 => "00011011",
 754 => "01111111",
 755 => "11110100",
 756 => "01011000",
 757 => "11000111",
 758 => "11101100",
 759 => "01101110",
 760 => "00011010",
 761 => "01011100",
 762 => "01011010",
 763 => "01100001",
 764 => "10111011",
 765 => "01000100",
 766 => "10011010",
 767 => "11100110",
 768 => "11100110",
 769 => "01110011",
 770 => "10100001",
 771 => "00010011",
 772 => "11001110",
 773 => "11000111",
 774 => "10001011",
 775 => "11010111",
 776 => "00111001",
 777 => "11011110",
 778 => "01110001",
 779 => "01111110",
 780 => "01100011",
 781 => "11010010",
 782 => "00100001",
 783 => "00111111",
 784 => "01010110",
 785 => "01110000",
 786 => "11110100",
 787 => "01011110",
 788 => "10000111",
 789 => "11101110",
 790 => "10101001",
 791 => "10100111",
 792 => "00111100",
 793 => "11010111",
 794 => "01001000",
 795 => "00010100",
 796 => "01111000",
 797 => "01000011",
 798 => "11000111",
 799 => "10111100",
 800 => "01000111",
 801 => "11011011",
 802 => "10001011",
 803 => "10011001",
 804 => "11010000",
 805 => "01100111",
 806 => "11000001",
 807 => "00101101",
 808 => "11000100",
 809 => "00011101",
 810 => "00011000",
 811 => "10010111",
 812 => "10010110",
 813 => "11001100",
 814 => "10100110",
 815 => "11110110",
 816 => "11100101",
 817 => "10000010",
 818 => "00011001",
 819 => "10111010",
 820 => "00010010",
 821 => "10111000",
 822 => "00011111",
 823 => "11011111",
 824 => "00001100",
 825 => "10001001",
 826 => "01000011",
 827 => "01110010",
 828 => "11000100",
 829 => "10100101",
 830 => "11111110",
 831 => "10011110",
 832 => "11110000",
 833 => "10010010",
 834 => "00001111",
 835 => "01010111",
 836 => "00110010",
 837 => "11011100",
 838 => "11000111",
 839 => "01011100",
 840 => "00001001",
 841 => "01100010",
 842 => "00100001",
 843 => "11010010",
 844 => "11100001",
 845 => "01100011",
 846 => "11000001",
 847 => "00000100",
 848 => "00110000",
 849 => "01100100",
 850 => "01010110",
 851 => "01110000",
 852 => "01110100",
 853 => "01000100",
 854 => "11100000",
 855 => "00000010",
 856 => "10000001",
 857 => "00111110",
 858 => "10000111",
 859 => "01110000",
 860 => "01010100",
 861 => "10010001",
 862 => "11001100",
 863 => "10011111",
 864 => "10111110",
 865 => "10100011",
 866 => "10110000",
 867 => "11100101",
 868 => "00100110",
 869 => "01111011",
 870 => "01111100",
 871 => "01100011",
 872 => "01010101",
 873 => "11000111",
 874 => "11001001",
 875 => "11000001",
 876 => "10111101",
 877 => "01111001",
 878 => "11101000",
 879 => "01000010",
 880 => "11100010",
 881 => "01000110",
 882 => "10011110",
 883 => "11101010",
 884 => "10111100",
 885 => "00100111",
 886 => "00110000",
 887 => "10011110",
 888 => "01110001",
 889 => "10101101",
 890 => "01000000",
 891 => "00000111",
 892 => "11101101",
 893 => "11101000",
 894 => "00110000",
 895 => "01111000",
 896 => "00111001",
 897 => "10000111",
 898 => "10111100",
 899 => "11011001",
 900 => "11000001",
 901 => "01101111",
 902 => "11101111",
 903 => "11010101",
 904 => "11010100",
 905 => "11001001",
 906 => "00001011",
 907 => "10011110",
 908 => "00000110",
 909 => "10101001",
 910 => "00000111",
 911 => "11110001",
 912 => "10100000",
 913 => "10001000",
 914 => "01000010",
 915 => "01000100",
 916 => "11111111",
 917 => "11100110",
 918 => "11000111",
 919 => "11101001",
 920 => "01111001",
 921 => "00101101",
 922 => "01001000",
 923 => "11000111",
 924 => "00111111",
 925 => "00110010",
 926 => "10001010",
 927 => "01101101",
 928 => "10011110",
 929 => "01110010",
 930 => "10011000",
 931 => "11101101",
 932 => "00100011",
 933 => "00111110",
 934 => "00010111",
 935 => "01101000",
 936 => "00010111",
 937 => "10001001",
 938 => "11011010",
 939 => "01111110",
 940 => "10001001",
 941 => "01100101",
 942 => "11011010",
 943 => "11111111",
 944 => "01110000",
 945 => "01000100",
 946 => "01011010",
 947 => "00011000",
 948 => "11101111",
 949 => "01101000",
 950 => "01111100",
 951 => "10110000",
 952 => "10111011",
 953 => "10111000",
 954 => "01000100",
 955 => "01001001",
 956 => "01111110",
 957 => "01100010",
 958 => "11100110",
 959 => "10101010",
 960 => "00100100",
 961 => "10010000",
 962 => "11010101",
 963 => "01010101",
 964 => "10110101",
 965 => "01000011",
 966 => "11011000",
 967 => "00110110",
 968 => "01000000",
 969 => "11110100",
 970 => "00011101",
 971 => "10110010",
 972 => "10110000",
 973 => "10111100",
 974 => "00011110",
 975 => "10000001",
 976 => "00110010",
 977 => "11011010",
 978 => "01100100",
 979 => "10100000",
 980 => "10111010",
 981 => "00010010",
 982 => "00011010",
 983 => "01001111",
 984 => "10101011",
 985 => "11011000",
 986 => "11010101",
 987 => "10101110",
 988 => "11111111",
 989 => "01001010",
 990 => "11011000",
 991 => "01000010",
 992 => "01000001",
 993 => "01100000",
 994 => "00011011",
 995 => "11010110",
 996 => "00100000",
 997 => "01010101",
 998 => "11100100",
 999 => "11010010",
 1000 => "00110100",
 1001 => "11111111",
 1002 => "01101001",
 1003 => "01000011",
 1004 => "10111111",
 1005 => "01100011",
 1006 => "01101111",
 1007 => "00100011",
 1008 => "11010001",
 1009 => "00011001",
 1010 => "10101111",
 1011 => "10001101",
 1012 => "00110011",
 1013 => "00001101",
 1014 => "00001001",
 1015 => "10111101",
 1016 => "01100111",
 1017 => "11111000",
 1018 => "10111010",
 1019 => "01110001",
 1020 => "11100111",
 1021 => "10000110",
 1022 => "11111100",
 1023 => "10010101",
 1024 => "01101100",
 1025 => "00110001",
 1026 => "00000100",
 1027 => "00111010",
 1028 => "11101100",
 1029 => "00100100",
 1030 => "00101010",
 1031 => "01100000",
 1032 => "00100010",
 1033 => "11010001",
 1034 => "10110100",
 1035 => "11111011",
 1036 => "01000110",
 1037 => "11001010",
 1038 => "11110100",
 1039 => "00001101",
 1040 => "11110011",
 1041 => "11010101",
 1042 => "10000100",
 1043 => "10111110",
 1044 => "11101000",
 1045 => "01101110",
 1046 => "10001101",
 1047 => "01000001",
 1048 => "10001001",
 1049 => "01001010",
 1050 => "01011000",
 1051 => "01001110",
 1052 => "11101001",
 1053 => "01110100",
 1054 => "00010001",
 1055 => "11101010",
 1056 => "01110011",
 1057 => "00011001",
 1058 => "11011111",
 1059 => "11111000",
 1060 => "00101100",
 1061 => "00010100",
 1062 => "10101010",
 1063 => "11110110",
 1064 => "00111110",
 1065 => "01111011",
 1066 => "01000000",
 1067 => "11011111",
 1068 => "00100101",
 1069 => "01001100",
 1070 => "01010001",
 1071 => "01000010",
 1072 => "10111101",
 1073 => "11111011",
 1074 => "00101001",
 1075 => "00100110",
 1076 => "01110011",
 1077 => "11100100",
 1078 => "01111101",
 1079 => "00011010",
 1080 => "00010111",
 1081 => "10010001",
 1082 => "11100111",
 1083 => "01000111",
 1084 => "10010000",
 1085 => "10000100",
 1086 => "01001000",
 1087 => "01000111",
 1088 => "00100101",
 1089 => "01101011",
 1090 => "01111010",
 1091 => "11111011",
 1092 => "11110011",
 1093 => "11101101",
 1094 => "10010111",
 1095 => "10110100",
 1096 => "10110010",
 1097 => "10001000",
 1098 => "11010111",
 1099 => "01101100",
 1100 => "00000010",
 1101 => "11110000",
 1102 => "01000011",
 1103 => "01010010",
 1104 => "01101010",
 1105 => "10111110",
 1106 => "11100110",
 1107 => "00110001",
 1108 => "11011101",
 1109 => "01001000",
 1110 => "00000111",
 1111 => "01101100",
 1112 => "10001100",
 1113 => "10010111",
 1114 => "10001010",
 1115 => "01000001",
 1116 => "01101101",
 1117 => "00111011",
 1118 => "10100111",
 1119 => "01011100",
 1120 => "10011000",
 1121 => "00010111",
 1122 => "11000110",
 1123 => "01100010",
 1124 => "11111001",
 1125 => "10100011",
 1126 => "10100001",
 1127 => "01110101",
 1128 => "00110101",
 1129 => "01001010",
 1130 => "10001101",
 1131 => "11010000",
 1132 => "10100100",
 1133 => "01011011",
 1134 => "01001000",
 1135 => "10010001",
 1136 => "11110101",
 1137 => "00111000",
 1138 => "10011010",
 1139 => "00111010",
 1140 => "01010111",
 1141 => "11111111",
 1142 => "00111111",
 1143 => "11000011",
 1144 => "00101000",
 1145 => "00101001",
 1146 => "11011011",
 1147 => "01110110",
 1148 => "00100001",
 1149 => "00000111",
 1150 => "00011110",
 1151 => "01010101",
 1152 => "01110111",
 1153 => "01101010",
 1154 => "11111111",
 1155 => "11001010",
 1156 => "10001011",
 1157 => "00011000",
 1158 => "00101101",
 1159 => "11100000",
 1160 => "00010100",
 1161 => "10101010",
 1162 => "00010000",
 1163 => "10101011",
 1164 => "10001110",
 1165 => "01001110",
 1166 => "11011001",
 1167 => "00111000",
 1168 => "11011110",
 1169 => "11100010",
 1170 => "10000111",
 1171 => "11101010",
 1172 => "01010100",
 1173 => "11110010",
 1174 => "01001111",
 1175 => "01000010",
 1176 => "01010001",
 1177 => "10100111",
 1178 => "01101101",
 1179 => "10011000",
 1180 => "01111110",
 1181 => "01010001",
 1182 => "10111111",
 1183 => "00100110",
 1184 => "10001111",
 1185 => "11000010",
 1186 => "10110011",
 1187 => "00110010",
 1188 => "01101010",
 1189 => "00111000",
 1190 => "00000011",
 1191 => "10010001",
 1192 => "01101111",
 1193 => "01001111",
 1194 => "00011110",
 1195 => "10110000",
 1196 => "11101111",
 1197 => "01110100",
 1198 => "11111110",
 1199 => "11000100",
 1200 => "11001010",
 1201 => "11100101",
 1202 => "01001011",
 1203 => "01001111",
 1204 => "01101011",
 1205 => "01111111",
 1206 => "11000010",
 1207 => "11101111",
 1208 => "11000011",
 1209 => "10110111",
 1210 => "01011111",
 1211 => "01101110",
 1212 => "00101101",
 1213 => "11100111",
 1214 => "01110101",
 1215 => "10000101",
 1216 => "00101010",
 1217 => "00110001",
 1218 => "01010001",
 1219 => "00100111",
 1220 => "11100001",
 1221 => "01110010",
 1222 => "10001011",
 1223 => "10110100",
 1224 => "00111100",
 1225 => "01000010",
 1226 => "11100000",
 1227 => "00110010",
 1228 => "01111100",
 1229 => "01101100",
 1230 => "11110010",
 1231 => "00110001",
 1232 => "00101100",
 1233 => "10101101",
 1234 => "01100101",
 1235 => "01001000",
 1236 => "01000111",
 1237 => "01011011",
 1238 => "00100000",
 1239 => "10000110",
 1240 => "11010101",
 1241 => "11011100",
 1242 => "00101101",
 1243 => "00001101",
 1244 => "10111101",
 1245 => "01111001",
 1246 => "10000000",
 1247 => "01011010",
 1248 => "10011110",
 1249 => "01010100",
 1250 => "11010001",
 1251 => "00011010",
 1252 => "01011010",
 1253 => "10111110",
 1254 => "10111110",
 1255 => "10011100",
 1256 => "01101111",
 1257 => "01101010",
 1258 => "01111110",
 1259 => "01111011",
 1260 => "11110001",
 1261 => "10010111",
 1262 => "11110011",
 1263 => "10110100",
 1264 => "10111000",
 1265 => "01001111",
 1266 => "00110110",
 1267 => "10010100",
 1268 => "01001110",
 1269 => "10010100",
 1270 => "10000110",
 1271 => "10011111",
 1272 => "00101110",
 1273 => "01001010",
 1274 => "11101110",
 1275 => "00101111",
 1276 => "01111101",
 1277 => "10000010",
 1278 => "10101011",
 1279 => "00111110",
 1280 => "11000101",
 1281 => "11111100",
 1282 => "00100010",
 1283 => "00111111",
 1284 => "11011001",
 1285 => "10011011",
 1286 => "01000010",
 1287 => "01011100",
 1288 => "01101010",
 1289 => "10101000",
 1290 => "00110110",
 1291 => "01011100",
 1292 => "10010100",
 1293 => "00010010",
 1294 => "10011001",
 1295 => "01010011",
 1296 => "00101100",
 1297 => "10010111",
 1298 => "00111001",
 1299 => "00101110",
 1300 => "01110110",
 1301 => "01111100",
 1302 => "11100110",
 1303 => "00101001",
 1304 => "00001000",
 1305 => "10110101",
 1306 => "00000100",
 1307 => "11111101",
 1308 => "01111011",
 1309 => "00110100",
 1310 => "00000101",
 1311 => "11111001",
 1312 => "00100110",
 1313 => "00011010",
 1314 => "01100000",
 1315 => "00111101",
 1316 => "10001111",
 1317 => "11111101",
 1318 => "10101011",
 1319 => "11011000",
 1320 => "11011101",
 1321 => "10000101",
 1322 => "10101000",
 1323 => "11010101",
 1324 => "00110101",
 1325 => "10111011",
 1326 => "01110110",
 1327 => "01011001",
 1328 => "01001011",
 1329 => "01100011",
 1330 => "10011000",
 1331 => "01011000",
 1332 => "10110111",
 1333 => "00010110",
 1334 => "00101110",
 1335 => "10100110",
 1336 => "10101101",
 1337 => "00000011",
 1338 => "00010011",
 1339 => "00010101",
 1340 => "01100111",
 1341 => "10110111",
 1342 => "10010000",
 1343 => "10011101",
 1344 => "11011010",
 1345 => "10000110",
 1346 => "00010000",
 1347 => "10101100",
 1348 => "10001011",
 1349 => "01001110",
 1350 => "11011010",
 1351 => "11011001",
 1352 => "01110010",
 1353 => "11110001",
 1354 => "01101111",
 1355 => "10000000",
 1356 => "11000001",
 1357 => "10100011",
 1358 => "00100110",
 1359 => "10110111",
 1360 => "10100000",
 1361 => "00101100",
 1362 => "01000011",
 1363 => "01111001",
 1364 => "01011010",
 1365 => "00011110",
 1366 => "00000001",
 1367 => "01100011",
 1368 => "10010100",
 1369 => "11000101",
 1370 => "01000101",
 1371 => "10110100",
 1372 => "10001100",
 1373 => "10101000",
 1374 => "00111011",
 1375 => "11000110",
 1376 => "11111110",
 1377 => "00001000",
 1378 => "01100000",
 1379 => "10111011",
 1380 => "10101111",
 1381 => "11000110",
 1382 => "10110001",
 1383 => "10100100",
 1384 => "01000110",
 1385 => "10001010",
 1386 => "00000100",
 1387 => "10100011",
 1388 => "00010000",
 1389 => "01010000",
 1390 => "00000111",
 1391 => "00111111",
 1392 => "00100001",
 1393 => "00001110",
 1394 => "11111100",
 1395 => "11000111",
 1396 => "01101000",
 1397 => "00111101",
 1398 => "10010001",
 1399 => "00111001",
 1400 => "00111010",
 1401 => "10000100",
 1402 => "01101010",
 1403 => "10110110",
 1404 => "01110010",
 1405 => "01100100",
 1406 => "10000111",
 1407 => "10101100",
 1408 => "00110001",
 1409 => "11111000",
 1410 => "00010100",
 1411 => "00110111",
 1412 => "10101111",
 1413 => "11010100",
 1414 => "10011001",
 1415 => "01001001",
 1416 => "00000101",
 1417 => "01000000",
 1418 => "01110000",
 1419 => "00001011",
 1420 => "01100011",
 1421 => "01010100",
 1422 => "00000000",
 1423 => "11010111",
 1424 => "11011101",
 1425 => "01110001",
 1426 => "01111001",
 1427 => "11000011",
 1428 => "11100111",
 1429 => "10000101",
 1430 => "11101100",
 1431 => "01000100",
 1432 => "00100011",
 1433 => "10011100",
 1434 => "10111001",
 1435 => "10001000",
 1436 => "11101100",
 1437 => "00011010",
 1438 => "11101101",
 1439 => "01000010",
 1440 => "00010000",
 1441 => "10101011",
 1442 => "11011011",
 1443 => "00001011",
 1444 => "10001000",
 1445 => "10100000",
 1446 => "11110011",
 1447 => "00101101",
 1448 => "11111101",
 1449 => "01110111",
 1450 => "00101101",
 1451 => "00011100",
 1452 => "10110101",
 1453 => "01110100",
 1454 => "10000010",
 1455 => "11111101",
 1456 => "10001100",
 1457 => "00100011",
 1458 => "11011101",
 1459 => "11001101",
 1460 => "00110001",
 1461 => "11110100",
 1462 => "11001100",
 1463 => "01100111",
 1464 => "01000000",
 1465 => "11010100",
 1466 => "11011110",
 1467 => "11100101",
 1468 => "11101111",
 1469 => "11110101",
 1470 => "10001110",
 1471 => "10110011",
 1472 => "11101100",
 1473 => "01100011",
 1474 => "01110111",
 1475 => "01110011",
 1476 => "10111100",
 1477 => "11001100",
 1478 => "01010100",
 1479 => "11001010",
 1480 => "01010011",
 1481 => "10010010",
 1482 => "10101101",
 1483 => "01000111",
 1484 => "00010111",
 1485 => "01100101",
 1486 => "00101010",
 1487 => "11111100",
 1488 => "11000101",
 1489 => "00101011",
 1490 => "10100001",
 1491 => "00011011",
 1492 => "00111111",
 1493 => "01100100",
 1494 => "10000001",
 1495 => "11011101",
 1496 => "11011100",
 1497 => "11001001",
 1498 => "10111101",
 1499 => "00101100",
 1500 => "11011100",
 1501 => "00001001",
 1502 => "10011001",
 1503 => "01010000",
 1504 => "10011100",
 1505 => "10010001",
 1506 => "01011111",
 1507 => "00100010",
 1508 => "11000111",
 1509 => "11111101",
 1510 => "01111010",
 1511 => "01000001",
 1512 => "10100110",
 1513 => "01001010",
 1514 => "10001100",
 1515 => "01100111",
 1516 => "01000011",
 1517 => "11110010",
 1518 => "10111000",
 1519 => "11010001",
 1520 => "01111001",
 1521 => "11100010",
 1522 => "10101000",
 1523 => "01100110",
 1524 => "00001101",
 1525 => "10010110",
 1526 => "00111100",
 1527 => "10110001",
 1528 => "00111010",
 1529 => "11011000",
 1530 => "11001011",
 1531 => "11100011",
 1532 => "10111100",
 1533 => "01011110",
 1534 => "11011100",
 1535 => "11011111",
 1536 => "01010011",
 1537 => "00011000",
 1538 => "11001100",
 1539 => "00100101",
 1540 => "10000100",
 1541 => "11001010",
 1542 => "10110101",
 1543 => "00001000",
 1544 => "11100001",
 1545 => "01010101",
 1546 => "10110011",
 1547 => "11100001",
 1548 => "10111110",
 1549 => "00011011",
 1550 => "11000100",
 1551 => "11000001",
 1552 => "01111011",
 1553 => "11010010",
 1554 => "10100111",
 1555 => "10000110",
 1556 => "00001100",
 1557 => "10100101",
 1558 => "01001011",
 1559 => "01111111",
 1560 => "01011111",
 1561 => "00100100",
 1562 => "01001110",
 1563 => "11011001",
 1564 => "11000101",
 1565 => "10101111",
 1566 => "10101101",
 1567 => "11011110",
 1568 => "01101010",
 1569 => "01110000",
 1570 => "01100100",
 1571 => "00000010",
 1572 => "11000101",
 1573 => "11010011",
 1574 => "01011011",
 1575 => "10100111",
 1576 => "10100110",
 1577 => "01010011",
 1578 => "00001101",
 1579 => "00101010",
 1580 => "10011001",
 1581 => "01011111",
 1582 => "01110110",
 1583 => "10001010",
 1584 => "11111011",
 1585 => "00010111",
 1586 => "01011111",
 1587 => "01101110",
 1588 => "10111010",
 1589 => "10010110",
 1590 => "11110000",
 1591 => "10000001",
 1592 => "11101101",
 1593 => "10011010",
 1594 => "00011010",
 1595 => "00100011",
 1596 => "11010001",
 1597 => "10011011",
 1598 => "11010011",
 1599 => "01100011",
 1600 => "01011101",
 1601 => "10010101",
 1602 => "11000010",
 1603 => "00111010",
 1604 => "00111011",
 1605 => "10001011",
 1606 => "00111100",
 1607 => "11001111",
 1608 => "11001111",
 1609 => "10011010",
 1610 => "01110010",
 1611 => "11010000",
 1612 => "01100011",
 1613 => "01101101",
 1614 => "10001011",
 1615 => "00101000",
 1616 => "10001110",
 1617 => "00001000",
 1618 => "11011000",
 1619 => "10100011",
 1620 => "11001000",
 1621 => "00010101",
 1622 => "10000100",
 1623 => "00001100",
 1624 => "01001011",
 1625 => "11000111",
 1626 => "10011100",
 1627 => "11111010",
 1628 => "00011011",
 1629 => "01000011",
 1630 => "11010010",
 1631 => "00001101",
 1632 => "10000001",
 1633 => "00011100",
 1634 => "00010110",
 1635 => "11111111",
 1636 => "01101010",
 1637 => "11111011",
 1638 => "10011001",
 1639 => "00001010",
 1640 => "00110100",
 1641 => "00010110",
 1642 => "01110111",
 1643 => "10100010",
 1644 => "11111010",
 1645 => "11111111",
 1646 => "10110110",
 1647 => "01011001",
 1648 => "01110100",
 1649 => "00110101",
 1650 => "10000111",
 1651 => "10000111",
 1652 => "11110010",
 1653 => "10001100",
 1654 => "11111110",
 1655 => "10001001",
 1656 => "11001111",
 1657 => "11111001",
 1658 => "11001010",
 1659 => "10000100",
 1660 => "10111010",
 1661 => "00000010",
 1662 => "01110011",
 1663 => "11000101",
 1664 => "11100010",
 1665 => "00110001",
 1666 => "01011100",
 1667 => "10000001",
 1668 => "10100101",
 1669 => "00111101",
 1670 => "00000011",
 1671 => "00010000",
 1672 => "11001111",
 1673 => "10100111",
 1674 => "11101101",
 1675 => "00110111",
 1676 => "10110111",
 1677 => "01101110",
 1678 => "11111111",
 1679 => "01000010",
 1680 => "10110101",
 1681 => "11100110",
 1682 => "10101101",
 1683 => "11001100",
 1684 => "11010010",
 1685 => "10110011",
 1686 => "11000011",
 1687 => "10101100",
 1688 => "10001000",
 1689 => "11100110",
 1690 => "00110111",
 1691 => "01110110",
 1692 => "01010101",
 1693 => "11111110",
 1694 => "10100110",
 1695 => "01111000",
 1696 => "01011001",
 1697 => "00100000",
 1698 => "00111001",
 1699 => "01100011",
 1700 => "00001111",
 1701 => "10111000",
 1702 => "00011100",
 1703 => "00101111",
 1704 => "10000010",
 1705 => "01110000",
 1706 => "01001111",
 1707 => "10110111",
 1708 => "11011110",
 1709 => "11101110",
 1710 => "10011101",
 1711 => "00001110",
 1712 => "11101100",
 1713 => "00111110",
 1714 => "10001101",
 1715 => "01001001",
 1716 => "11101111",
 1717 => "10100100",
 1718 => "01010111",
 1719 => "11010110",
 1720 => "10000101",
 1721 => "11001000",
 1722 => "01001101",
 1723 => "00001000",
 1724 => "11100011",
 1725 => "10101011",
 1726 => "00001010",
 1727 => "10111110",
 1728 => "11110111",
 1729 => "00001111",
 1730 => "00011000",
 1731 => "10110100",
 1732 => "10000011",
 1733 => "11010001",
 1734 => "01111110",
 1735 => "10101011",
 1736 => "01100110",
 1737 => "01111101",
 1738 => "01101110",
 1739 => "11110101",
 1740 => "11010110",
 1741 => "10010001",
 1742 => "00101011",
 1743 => "10101010",
 1744 => "11011111",
 1745 => "11110111",
 1746 => "10000001",
 1747 => "11000001",
 1748 => "10111010",
 1749 => "11000000",
 1750 => "00000111",
 1751 => "11001101",
 1752 => "00000101",
 1753 => "10011011",
 1754 => "01011110",
 1755 => "10011011",
 1756 => "00000101",
 1757 => "00111011",
 1758 => "11100011",
 1759 => "11111011",
 1760 => "10010011",
 1761 => "00110000",
 1762 => "00010110",
 1763 => "01011100",
 1764 => "11111011",
 1765 => "10001010",
 1766 => "10110010",
 1767 => "00110011",
 1768 => "01110000",
 1769 => "10010100",
 1770 => "11111100",
 1771 => "00101110",
 1772 => "10001111",
 1773 => "00011010",
 1774 => "11010011",
 1775 => "10001011",
 1776 => "00101110",
 1777 => "00010010",
 1778 => "00011110",
 1779 => "01100110",
 1780 => "10000110",
 1781 => "00110111",
 1782 => "10011001",
 1783 => "00110000",
 1784 => "10001000",
 1785 => "00100011",
 1786 => "11101011",
 1787 => "11110011",
 1788 => "00110010",
 1789 => "10101000",
 1790 => "10011110",
 1791 => "11111100",
 1792 => "10001010",
 1793 => "10110101",
 1794 => "01101101",
 1795 => "11010011",
 1796 => "10101110",
 1797 => "10010011",
 1798 => "01001101",
 1799 => "00111101",
 1800 => "10010111",
 1801 => "11000110",
 1802 => "00111111",
 1803 => "10100110",
 1804 => "10111100",
 1805 => "10010011",
 1806 => "00101010",
 1807 => "10001100",
 1808 => "10011110",
 1809 => "01000011",
 1810 => "10110100",
 1811 => "10010111",
 1812 => "01100100",
 1813 => "11110011",
 1814 => "11010001",
 1815 => "11100000",
 1816 => "01001100",
 1817 => "01001100",
 1818 => "00001001",
 1819 => "01100100",
 1820 => "10001001",
 1821 => "01001000",
 1822 => "10001010",
 1823 => "11101100",
 1824 => "11001100",
 1825 => "00111100",
 1826 => "10011001",
 1827 => "10101100",
 1828 => "11000101",
 1829 => "11110001",
 1830 => "10100011",
 1831 => "01111101",
 1832 => "10110100",
 1833 => "11111011",
 1834 => "00001111",
 1835 => "01001011",
 1836 => "01000101",
 1837 => "10100111",
 1838 => "01000111",
 1839 => "00000101",
 1840 => "11000100",
 1841 => "10110010",
 1842 => "00011010",
 1843 => "01001001",
 1844 => "01011100",
 1845 => "11000100",
 1846 => "11000101",
 1847 => "10101000",
 1848 => "00110000",
 1849 => "01001100",
 1850 => "01100100",
 1851 => "01111100",
 1852 => "10011011",
 1853 => "11011000",
 1854 => "00010111",
 1855 => "00000000",
 1856 => "00100001",
 1857 => "00110000",
 1858 => "10000101",
 1859 => "10100110",
 1860 => "11111010",
 1861 => "01011000",
 1862 => "11111000",
 1863 => "10110011",
 1864 => "00010010",
 1865 => "11100011",
 1866 => "10000001",
 1867 => "00110011",
 1868 => "11010001",
 1869 => "01100111",
 1870 => "11011111",
 1871 => "10101111",
 1872 => "00001101",
 1873 => "10110101",
 1874 => "00011110",
 1875 => "01101101",
 1876 => "11000011",
 1877 => "00100111",
 1878 => "01100010",
 1879 => "01111010",
 1880 => "01000000",
 1881 => "00011000",
 1882 => "01101111",
 1883 => "00101101",
 1884 => "00000010",
 1885 => "10010101",
 1886 => "10100011",
 1887 => "01010101",
 1888 => "01011111",
 1889 => "00111111",
 1890 => "01100000",
 1891 => "11001111",
 1892 => "11001100",
 1893 => "11100111",
 1894 => "11110100",
 1895 => "01011010",
 1896 => "01110101",
 1897 => "00001011",
 1898 => "11110101",
 1899 => "10101111",
 1900 => "10000101",
 1901 => "00101110",
 1902 => "00110000",
 1903 => "11100000",
 1904 => "01000010",
 1905 => "00111100",
 1906 => "00001100",
 1907 => "10011010",
 1908 => "10100000",
 1909 => "01010101",
 1910 => "00010001",
 1911 => "01010101",
 1912 => "01111101",
 1913 => "00110101",
 1914 => "01111011",
 1915 => "00110011",
 1916 => "00011110",
 1917 => "10001010",
 1918 => "11100000",
 1919 => "10001101",
 1920 => "11101111",
 1921 => "10011011",
 1922 => "10110111",
 1923 => "10100101",
 1924 => "01101101",
 1925 => "01011000",
 1926 => "10010100",
 1927 => "01101101",
 1928 => "00111011",
 1929 => "01010101",
 1930 => "11001111",
 1931 => "11010100",
 1932 => "01010111",
 1933 => "10010111",
 1934 => "11001010",
 1935 => "10111111",
 1936 => "10001010",
 1937 => "01000011",
 1938 => "01100110",
 1939 => "00100000",
 1940 => "01110010",
 1941 => "10101000",
 1942 => "11111001",
 1943 => "00010100",
 1944 => "10001001",
 1945 => "01010101",
 1946 => "00111001",
 1947 => "00011110",
 1948 => "01000111",
 1949 => "01111001",
 1950 => "00101010",
 1951 => "01011011",
 1952 => "11011010",
 1953 => "00010000",
 1954 => "01010110",
 1955 => "01001100",
 1956 => "10011111",
 1957 => "10100010",
 1958 => "01001000",
 1959 => "00010110",
 1960 => "00101100",
 1961 => "10111010",
 1962 => "10110100",
 1963 => "11010010",
 1964 => "00110000",
 1965 => "00011111",
 1966 => "10001011",
 1967 => "01111000",
 1968 => "01010111",
 1969 => "11111110",
 1970 => "01101111",
 1971 => "10000011",
 1972 => "10010010",
 1973 => "00101111",
 1974 => "00101100",
 1975 => "01000000",
 1976 => "11000001",
 1977 => "11100001",
 1978 => "01010111",
 1979 => "11100011",
 1980 => "01011110",
 1981 => "11101110",
 1982 => "11000100",
 1983 => "11001010",
 1984 => "10101001",
 1985 => "00110000",
 1986 => "10101010",
 1987 => "00010011",
 1988 => "10000001",
 1989 => "00110010",
 1990 => "10011000",
 1991 => "10100001",
 1992 => "11111100",
 1993 => "01011110",
 1994 => "01000111",
 1995 => "10111110",
 1996 => "00111110",
 1997 => "01100000",
 1998 => "01111000",
 1999 => "10111111",
 2000 => "10110101",
 2001 => "11111010",
 2002 => "11101011",
 2003 => "01010011",
 2004 => "10111100",
 2005 => "01100000",
 2006 => "10111110",
 2007 => "10111000",
 2008 => "11010000",
 2009 => "11011010",
 2010 => "01011110",
 2011 => "11001010",
 2012 => "00100011",
 2013 => "10011001",
 2014 => "11101011",
 2015 => "11001000",
 2016 => "11100000",
 2017 => "10011011",
 2018 => "11111100",
 2019 => "00001001",
 2020 => "11011011",
 2021 => "00001000",
 2022 => "11000101",
 2023 => "01011111",
 2024 => "10000001",
 2025 => "00010111",
 2026 => "10110111",
 2027 => "10001100",
 2028 => "00110110",
 2029 => "10011100",
 2030 => "00000100",
 2031 => "10011111",
 2032 => "10010100",
 2033 => "00110101",
 2034 => "11110101",
 2035 => "01100111",
 2036 => "10001001",
 2037 => "11101000",
 2038 => "01000100",
 2039 => "10100000",
 2040 => "00010101",
 2041 => "01100100",
 2042 => "11001011",
 2043 => "00000100",
 2044 => "10101001",
 2045 => "00001001",
 2046 => "00011110",
 2047 => "01111100",
 2048 => "00011001",
 2049 => "00000001",
 2050 => "00110000",
 2051 => "01010100",
 2052 => "00111000",
 2053 => "11110111",
 2054 => "11010011",
 2055 => "00100111",
 2056 => "10111100",
 2057 => "01011110",
 2058 => "10000010",
 2059 => "01110110",
 2060 => "10010000",
 2061 => "00111111",
 2062 => "01001100",
 2063 => "11100010",
 2064 => "01100100",
 2065 => "00101110",
 2066 => "10011110",
 2067 => "01000010",
 2068 => "11100001",
 2069 => "11001010",
 2070 => "01111001",
 2071 => "11000010",
 2072 => "01101111",
 2073 => "01011100",
 2074 => "11100010",
 2075 => "11011010",
 2076 => "00111011",
 2077 => "00110111",
 2078 => "01010010",
 2079 => "01111100",
 2080 => "00100010",
 2081 => "10101110",
 2082 => "11100000",
 2083 => "01110010",
 2084 => "11110000",
 2085 => "01101100",
 2086 => "10000000",
 2087 => "11000011",
 2088 => "01100101",
 2089 => "00110011",
 2090 => "10010110",
 2091 => "00110101",
 2092 => "11011001",
 2093 => "11110100",
 2094 => "11101110",
 2095 => "11111110",
 2096 => "11110101",
 2097 => "11001001",
 2098 => "10111011",
 2099 => "01110010",
 2100 => "01011101",
 2101 => "00100111",
 2102 => "10010110",
 2103 => "00110111",
 2104 => "10011001",
 2105 => "01111101",
 2106 => "11010000",
 2107 => "00001001",
 2108 => "10110100",
 2109 => "11011000",
 2110 => "00001011",
 2111 => "01111000",
 2112 => "00010001",
 2113 => "11010100",
 2114 => "00000110",
 2115 => "01100000",
 2116 => "10011011",
 2117 => "11110100",
 2118 => "10101101",
 2119 => "00101011",
 2120 => "01110001",
 2121 => "10011110",
 2122 => "00011000",
 2123 => "11000110",
 2124 => "01010110",
 2125 => "01111100",
 2126 => "10110101",
 2127 => "10111101",
 2128 => "11011000",
 2129 => "00100100",
 2130 => "00110001",
 2131 => "10010100",
 2132 => "01100111",
 2133 => "01100111",
 2134 => "01100011",
 2135 => "10101001",
 2136 => "01100000",
 2137 => "10111010",
 2138 => "11101000",
 2139 => "11101001",
 2140 => "10100101",
 2141 => "00101011",
 2142 => "01010110",
 2143 => "00100111",
 2144 => "00100011",
 2145 => "01111101",
 2146 => "00011101",
 2147 => "10111000",
 2148 => "01001100",
 2149 => "11100101",
 2150 => "10111100",
 2151 => "01010000",
 2152 => "11010011",
 2153 => "10010001",
 2154 => "10110010",
 2155 => "00100010",
 2156 => "10000001",
 2157 => "00010000",
 2158 => "10000011",
 2159 => "00001011",
 2160 => "11010111",
 2161 => "10100010",
 2162 => "11010110",
 2163 => "01111100",
 2164 => "01011010",
 2165 => "01111001",
 2166 => "10011110",
 2167 => "10111010",
 2168 => "10010000",
 2169 => "11010001",
 2170 => "11000101",
 2171 => "00001001",
 2172 => "01001010",
 2173 => "10000001",
 2174 => "11100100",
 2175 => "01010001",
 2176 => "10101111",
 2177 => "11010100",
 2178 => "01001110",
 2179 => "11001111",
 2180 => "11110001",
 2181 => "10010000",
 2182 => "01110011",
 2183 => "01101101",
 2184 => "00010000",
 2185 => "01011010",
 2186 => "11111111",
 2187 => "11101001",
 2188 => "01000101",
 2189 => "11100000",
 2190 => "01010001",
 2191 => "10101010",
 2192 => "01011011",
 2193 => "00101110",
 2194 => "01110111",
 2195 => "00100010",
 2196 => "01000110",
 2197 => "10111001",
 2198 => "01110100",
 2199 => "11100011",
 2200 => "01100111",
 2201 => "00101000",
 2202 => "01000101",
 2203 => "10101111",
 2204 => "11110011",
 2205 => "00010110",
 2206 => "11100000",
 2207 => "01010011",
 2208 => "11001111",
 2209 => "11101001",
 2210 => "01111101",
 2211 => "11010110",
 2212 => "10100001",
 2213 => "01111110",
 2214 => "01010101",
 2215 => "10101010",
 2216 => "00010110",
 2217 => "11000000",
 2218 => "00011010",
 2219 => "11010000",
 2220 => "10011000",
 2221 => "01001000",
 2222 => "00000100",
 2223 => "10010011",
 2224 => "10100110",
 2225 => "11111010",
 2226 => "00100110",
 2227 => "11000111",
 2228 => "10101010",
 2229 => "11011110",
 2230 => "00000001",
 2231 => "11011101",
 2232 => "00000011",
 2233 => "01100010",
 2234 => "00101111",
 2235 => "11001110",
 2236 => "11001010",
 2237 => "01000101",
 2238 => "10110010",
 2239 => "10011100",
 2240 => "00110101",
 2241 => "01110010",
 2242 => "00010001",
 2243 => "01110100",
 2244 => "01000111",
 2245 => "01001011",
 2246 => "10001100",
 2247 => "11101011",
 2248 => "01101011",
 2249 => "00011111",
 2250 => "11101101",
 2251 => "11001010",
 2252 => "01111110",
 2253 => "11001010",
 2254 => "11011111",
 2255 => "01011110",
 2256 => "10101111",
 2257 => "01000110",
 2258 => "01101010",
 2259 => "00000101",
 2260 => "01000100",
 2261 => "01110110",
 2262 => "11101110",
 2263 => "01100000",
 2264 => "11011000",
 2265 => "01010110",
 2266 => "01100101",
 2267 => "00110101",
 2268 => "00000111",
 2269 => "11010000",
 2270 => "01000011",
 2271 => "00010001",
 2272 => "10000000",
 2273 => "01110101",
 2274 => "11100110",
 2275 => "00100110",
 2276 => "01110001",
 2277 => "01100111",
 2278 => "10110011",
 2279 => "01001110",
 2280 => "11111100",
 2281 => "01011100",
 2282 => "01001001",
 2283 => "11100110",
 2284 => "10000010",
 2285 => "10001111",
 2286 => "11010001",
 2287 => "11101110",
 2288 => "10000101",
 2289 => "00110010",
 2290 => "01101110",
 2291 => "10110111",
 2292 => "01011011",
 2293 => "10111000",
 2294 => "10101101",
 2295 => "10110111",
 2296 => "11001001",
 2297 => "00101110",
 2298 => "11110000",
 2299 => "01000000",
 2300 => "11011010",
 2301 => "11100011",
 2302 => "01101001",
 2303 => "01011101",
 2304 => "00110010",
 2305 => "01001101",
 2306 => "10100001",
 2307 => "01001110",
 2308 => "11101101",
 2309 => "00000000",
 2310 => "00101111",
 2311 => "10010111",
 2312 => "00110111",
 2313 => "11001011",
 2314 => "00001100",
 2315 => "00000010",
 2316 => "01000000",
 2317 => "01001111",
 2318 => "00110111",
 2319 => "10110100",
 2320 => "10001110",
 2321 => "11010101",
 2322 => "01111011",
 2323 => "11010001",
 2324 => "01000010",
 2325 => "00100001",
 2326 => "01100010",
 2327 => "01011111",
 2328 => "00100100",
 2329 => "00100100",
 2330 => "11010100",
 2331 => "11010001",
 2332 => "11001111",
 2333 => "10010110",
 2334 => "11011111",
 2335 => "01001110",
 2336 => "10011000",
 2337 => "00101000",
 2338 => "01100011",
 2339 => "00111101",
 2340 => "00111111",
 2341 => "11011101",
 2342 => "00110011",
 2343 => "00110010",
 2344 => "10001000",
 2345 => "00011101",
 2346 => "01101001",
 2347 => "10001011",
 2348 => "00100010",
 2349 => "10000010",
 2350 => "01000000",
 2351 => "01110111",
 2352 => "00010111",
 2353 => "10010000",
 2354 => "00101100",
 2355 => "01111001",
 2356 => "00111001",
 2357 => "00101100",
 2358 => "11010111",
 2359 => "10100000",
 2360 => "11000100",
 2361 => "10001000",
 2362 => "01001110",
 2363 => "10011010",
 2364 => "01101100",
 2365 => "11011111",
 2366 => "10111101",
 2367 => "10001000",
 2368 => "10100110",
 2369 => "10110000",
 2370 => "00111011",
 2371 => "01001000",
 2372 => "00100101",
 2373 => "00000010",
 2374 => "10000011",
 2375 => "00010000",
 2376 => "01000111",
 2377 => "10001110",
 2378 => "11100010",
 2379 => "00001101",
 2380 => "10100010",
 2381 => "10001110",
 2382 => "11110000",
 2383 => "10011000",
 2384 => "01111110",
 2385 => "10010011",
 2386 => "00011111",
 2387 => "00100010",
 2388 => "11100001",
 2389 => "01100110",
 2390 => "01101101",
 2391 => "00110001",
 2392 => "01111110",
 2393 => "10101100",
 2394 => "00011000",
 2395 => "00001110",
 2396 => "00011110",
 2397 => "00101000",
 2398 => "10110101",
 2399 => "00100111",
 2400 => "01001111",
 2401 => "01001001",
 2402 => "11111101",
 2403 => "10111011",
 2404 => "01111111",
 2405 => "10101001",
 2406 => "00001010",
 2407 => "10011001",
 2408 => "01100000",
 2409 => "00100001",
 2410 => "11001011",
 2411 => "00001001",
 2412 => "01011100",
 2413 => "01001001",
 2414 => "11001100",
 2415 => "00111010",
 2416 => "11000001",
 2417 => "00100100",
 2418 => "00110110",
 2419 => "11100111",
 2420 => "11001101",
 2421 => "00001001",
 2422 => "00101000",
 2423 => "11100011",
 2424 => "10000011",
 2425 => "11001111",
 2426 => "11100010",
 2427 => "01101101",
 2428 => "01100000",
 2429 => "01010110",
 2430 => "00101000",
 2431 => "10001101",
 2432 => "10100111",
 2433 => "11010011",
 2434 => "01011101",
 2435 => "01010101",
 2436 => "11001000",
 2437 => "00101001",
 2438 => "01110111",
 2439 => "10011110",
 2440 => "10000111",
 2441 => "00001010",
 2442 => "01111111",
 2443 => "00111100",
 2444 => "10001001",
 2445 => "00011000",
 2446 => "01000110",
 2447 => "11001000",
 2448 => "00000101",
 2449 => "11011111",
 2450 => "10100001",
 2451 => "10100000",
 2452 => "10101010",
 2453 => "01110110",
 2454 => "00100001",
 2455 => "00010110",
 2456 => "00001100",
 2457 => "00010000",
 2458 => "01111010",
 2459 => "00001101",
 2460 => "00000010",
 2461 => "10000100",
 2462 => "11001110",
 2463 => "00110010",
 2464 => "11010001",
 2465 => "11010111",
 2466 => "01101000",
 2467 => "11000010",
 2468 => "00100111",
 2469 => "11010110",
 2470 => "11001011",
 2471 => "11010001",
 2472 => "10000000",
 2473 => "11111110",
 2474 => "11010101",
 2475 => "10101110",
 2476 => "00011101",
 2477 => "10110100",
 2478 => "01010111",
 2479 => "11111001",
 2480 => "00011010",
 2481 => "01011001",
 2482 => "01101101",
 2483 => "00000111",
 2484 => "01111111",
 2485 => "01110111",
 2486 => "00001111",
 2487 => "11100011",
 2488 => "00000010",
 2489 => "10000000",
 2490 => "11111000",
 2491 => "00011100",
 2492 => "10100011",
 2493 => "00101011",
 2494 => "01010110",
 2495 => "10100111",
 2496 => "10100100",
 2497 => "00011110",
 2498 => "10111101",
 2499 => "00101011",
 2500 => "00111010",
 2501 => "01010110",
 2502 => "11011011",
 2503 => "10011111",
 2504 => "10011010",
 2505 => "00010011",
 2506 => "11001010",
 2507 => "00001111",
 2508 => "10111001",
 2509 => "01101111",
 2510 => "11101111",
 2511 => "00100010",
 2512 => "00011010",
 2513 => "11110000",
 2514 => "11010101",
 2515 => "11010000",
 2516 => "00001110",
 2517 => "11011110",
 2518 => "11100011",
 2519 => "01011010",
 2520 => "00111001",
 2521 => "11011111",
 2522 => "10000011",
 2523 => "10010011",
 2524 => "01101100",
 2525 => "00100110",
 2526 => "01101100",
 2527 => "00001111",
 2528 => "00111010",
 2529 => "11110011",
 2530 => "10110101",
 2531 => "10010101",
 2532 => "11110010",
 2533 => "01110010",
 2534 => "01011101",
 2535 => "10001011",
 2536 => "00110111",
 2537 => "11000111",
 2538 => "11101111",
 2539 => "01011101",
 2540 => "10101101",
 2541 => "11001001",
 2542 => "01100011",
 2543 => "11110110",
 2544 => "00100010",
 2545 => "10101011",
 2546 => "01111111",
 2547 => "01001111",
 2548 => "10101011",
 2549 => "01111111",
 2550 => "01100101",
 2551 => "11000010",
 2552 => "11000101",
 2553 => "01000001",
 2554 => "10001011",
 2555 => "01001010",
 2556 => "01100110",
 2557 => "01011010",
 2558 => "00011111",
 2559 => "10110000",
 2560 => "11010011",
 2561 => "01001101",
 2562 => "01111100",
 2563 => "11000001",
 2564 => "00000101",
 2565 => "01010011",
 2566 => "11011110",
 2567 => "11111100",
 2568 => "00101001",
 2569 => "11111111",
 2570 => "10111001",
 2571 => "01011001",
 2572 => "01110011",
 2573 => "01100101",
 2574 => "11001101",
 2575 => "00010000",
 2576 => "00100001",
 2577 => "11110110",
 2578 => "11010111",
 2579 => "00011001",
 2580 => "11101101",
 2581 => "10011010",
 2582 => "01010011",
 2583 => "00111000",
 2584 => "10000101",
 2585 => "10111011",
 2586 => "10100011",
 2587 => "10000010",
 2588 => "00000101",
 2589 => "01101101",
 2590 => "00011001",
 2591 => "10010000",
 2592 => "10110101",
 2593 => "10001011",
 2594 => "10011110",
 2595 => "11100000",
 2596 => "00001000",
 2597 => "01001001",
 2598 => "01101010",
 2599 => "10010010",
 2600 => "10001111",
 2601 => "00111110",
 2602 => "11110010",
 2603 => "00001100",
 2604 => "10010111",
 2605 => "11111001",
 2606 => "00001010",
 2607 => "01110010",
 2608 => "01100001",
 2609 => "10010001",
 2610 => "11110110",
 2611 => "01101101",
 2612 => "01101010",
 2613 => "10011011",
 2614 => "01010110",
 2615 => "00101010",
 2616 => "01100110",
 2617 => "01010011",
 2618 => "00010101",
 2619 => "11011011",
 2620 => "01101001",
 2621 => "00110011",
 2622 => "01001011",
 2623 => "01001001",
 2624 => "00110000",
 2625 => "01101101",
 2626 => "01111111",
 2627 => "01100001",
 2628 => "10010010",
 2629 => "11100011",
 2630 => "11111010",
 2631 => "01010111",
 2632 => "11010010",
 2633 => "10010101",
 2634 => "01100001",
 2635 => "11001101",
 2636 => "01111001",
 2637 => "10010111",
 2638 => "11111100",
 2639 => "10111110",
 2640 => "01001000",
 2641 => "11110010",
 2642 => "00100010",
 2643 => "10101110",
 2644 => "11101000",
 2645 => "01100100",
 2646 => "10001110",
 2647 => "00110000",
 2648 => "10101111",
 2649 => "11011100",
 2650 => "01110010",
 2651 => "10011001",
 2652 => "10111111",
 2653 => "00010100",
 2654 => "11111001",
 2655 => "10011110",
 2656 => "10101010",
 2657 => "01101111",
 2658 => "10110001",
 2659 => "10010110",
 2660 => "00001111",
 2661 => "11111001",
 2662 => "01100011",
 2663 => "00000001",
 2664 => "00100110",
 2665 => "11001101",
 2666 => "10000001",
 2667 => "01111111",
 2668 => "10111001",
 2669 => "11101001",
 2670 => "01101110",
 2671 => "00101111",
 2672 => "10001110",
 2673 => "10111100",
 2674 => "10000111",
 2675 => "00010101",
 2676 => "00000111",
 2677 => "00001001",
 2678 => "00110100",
 2679 => "01010101",
 2680 => "01111101",
 2681 => "00011001",
 2682 => "11001100",
 2683 => "11101111",
 2684 => "00110111",
 2685 => "01011000",
 2686 => "00101110",
 2687 => "10011101",
 2688 => "00010000",
 2689 => "00110110",
 2690 => "00100111",
 2691 => "01011010",
 2692 => "11011000",
 2693 => "01111001",
 2694 => "11010110",
 2695 => "00101000",
 2696 => "10011010",
 2697 => "00001101",
 2698 => "10110100",
 2699 => "00100111",
 2700 => "11001111",
 2701 => "11011101",
 2702 => "10011111",
 2703 => "01101100",
 2704 => "10001011",
 2705 => "00010000",
 2706 => "11011000",
 2707 => "10101111",
 2708 => "00100110",
 2709 => "10010010",
 2710 => "00101011",
 2711 => "00100010",
 2712 => "10001111",
 2713 => "01011110",
 2714 => "11110011",
 2715 => "00100001",
 2716 => "11100010",
 2717 => "00000011",
 2718 => "00001011",
 2719 => "01100001",
 2720 => "10100000",
 2721 => "01000000",
 2722 => "01111001",
 2723 => "11011001",
 2724 => "01101100",
 2725 => "01110010",
 2726 => "01001001",
 2727 => "10010001",
 2728 => "01011101",
 2729 => "10111010",
 2730 => "01101101",
 2731 => "10111101",
 2732 => "00100010",
 2733 => "01011000",
 2734 => "10100001",
 2735 => "10100001",
 2736 => "00000100",
 2737 => "10010010",
 2738 => "01111101",
 2739 => "11101101",
 2740 => "10110111",
 2741 => "11001101",
 2742 => "00111111",
 2743 => "10100111",
 2744 => "10101110",
 2745 => "10001110",
 2746 => "10000011",
 2747 => "10011001",
 2748 => "10010111",
 2749 => "11100010",
 2750 => "11100000",
 2751 => "11001111",
 2752 => "10101101",
 2753 => "10101010",
 2754 => "10100111",
 2755 => "11000110",
 2756 => "10010110",
 2757 => "10110011",
 2758 => "00011101",
 2759 => "01110011",
 2760 => "10100110",
 2761 => "00011110",
 2762 => "10010110",
 2763 => "10011011",
 2764 => "10111010",
 2765 => "01001000",
 2766 => "00101001",
 2767 => "11000001",
 2768 => "01001110",
 2769 => "01110011",
 2770 => "00100011",
 2771 => "01000001",
 2772 => "10000000",
 2773 => "10100100",
 2774 => "00111001",
 2775 => "01010000",
 2776 => "11101101",
 2777 => "01011001",
 2778 => "00110011",
 2779 => "00111101",
 2780 => "00101111",
 2781 => "00001001",
 2782 => "11111111",
 2783 => "11001000",
 2784 => "01111111",
 2785 => "10100000",
 2786 => "10000011",
 2787 => "00110000",
 2788 => "00001100",
 2789 => "11000111",
 2790 => "01000100",
 2791 => "01110101",
 2792 => "00011001",
 2793 => "11100010",
 2794 => "00111101",
 2795 => "10111110",
 2796 => "11011100",
 2797 => "10000011",
 2798 => "10001011",
 2799 => "11111101",
 2800 => "01011100",
 2801 => "11111100",
 2802 => "00011110",
 2803 => "01011011",
 2804 => "01100110",
 2805 => "11110100",
 2806 => "11011000",
 2807 => "10000010",
 2808 => "00111110",
 2809 => "00011001",
 2810 => "11010011",
 2811 => "10010000",
 2812 => "11110111",
 2813 => "11111001",
 2814 => "11101011",
 2815 => "00000011",
 2816 => "01101011",
 2817 => "11010001",
 2818 => "11000001",
 2819 => "01101011",
 2820 => "00001111",
 2821 => "01011101",
 2822 => "01100001",
 2823 => "10010010",
 2824 => "11001110",
 2825 => "10101001",
 2826 => "01100011",
 2827 => "10110100",
 2828 => "00010010",
 2829 => "11110110",
 2830 => "00110111",
 2831 => "11101011",
 2832 => "11011110",
 2833 => "10100011",
 2834 => "00111010",
 2835 => "00010100",
 2836 => "00110000",
 2837 => "10100011",
 2838 => "11110101",
 2839 => "11011010",
 2840 => "00000110",
 2841 => "11111000",
 2842 => "01110101",
 2843 => "00001000",
 2844 => "10110101",
 2845 => "11111001",
 2846 => "11010101",
 2847 => "01100011",
 2848 => "01011111",
 2849 => "01110011",
 2850 => "00011111",
 2851 => "00100000",
 2852 => "00001010",
 2853 => "10000000",
 2854 => "00001100",
 2855 => "01111011",
 2856 => "11101110",
 2857 => "11100000",
 2858 => "10011011",
 2859 => "10001000",
 2860 => "00110101",
 2861 => "00010101",
 2862 => "11010001",
 2863 => "10110000",
 2864 => "01110010",
 2865 => "00000101",
 2866 => "10101110",
 2867 => "10010010",
 2868 => "01100000",
 2869 => "10100011",
 2870 => "01111111",
 2871 => "10110010",
 2872 => "11110000",
 2873 => "01110101",
 2874 => "11000011",
 2875 => "01100100",
 2876 => "11100110",
 2877 => "00000011",
 2878 => "10100101",
 2879 => "11010010",
 2880 => "01101000",
 2881 => "10001000",
 2882 => "10110111",
 2883 => "01010110",
 2884 => "01111011",
 2885 => "00011000",
 2886 => "01001001",
 2887 => "00000110",
 2888 => "01101111",
 2889 => "01001111",
 2890 => "01001010",
 2891 => "00101111",
 2892 => "01000000",
 2893 => "00101110",
 2894 => "00110000",
 2895 => "00010101",
 2896 => "00000110",
 2897 => "00100011",
 2898 => "01101011",
 2899 => "11110010",
 2900 => "00111001",
 2901 => "10100011",
 2902 => "10000101",
 2903 => "01101010",
 2904 => "10110111",
 2905 => "11110010",
 2906 => "01111000",
 2907 => "11001001",
 2908 => "10001110",
 2909 => "10001101",
 2910 => "01011101",
 2911 => "00100101",
 2912 => "00110001",
 2913 => "11110110",
 2914 => "00101100",
 2915 => "11010111",
 2916 => "11010001",
 2917 => "11110101",
 2918 => "11101011",
 2919 => "00110111",
 2920 => "01000000",
 2921 => "01011101",
 2922 => "10100111",
 2923 => "00100011",
 2924 => "01010101",
 2925 => "11100100",
 2926 => "10011011",
 2927 => "00011001",
 2928 => "10100001",
 2929 => "00001001",
 2930 => "01110100",
 2931 => "00001100",
 2932 => "01110110",
 2933 => "10101011",
 2934 => "00110011",
 2935 => "01100100",
 2936 => "11110011",
 2937 => "11010010",
 2938 => "01001101",
 2939 => "10011101",
 2940 => "01011010",
 2941 => "00010001",
 2942 => "01111100",
 2943 => "10011101",
 2944 => "11100000",
 2945 => "10110111",
 2946 => "00101110",
 2947 => "10110110",
 2948 => "10010100",
 2949 => "11111100",
 2950 => "11011001",
 2951 => "11111110",
 2952 => "00000000",
 2953 => "11011001",
 2954 => "10100011",
 2955 => "00100111",
 2956 => "10110111",
 2957 => "10101100",
 2958 => "10000011",
 2959 => "01111001",
 2960 => "01110000",
 2961 => "01111010",
 2962 => "01100110",
 2963 => "10010011",
 2964 => "01100100",
 2965 => "01100100",
 2966 => "00011011",
 2967 => "00010101",
 2968 => "01011111",
 2969 => "01001011",
 2970 => "11100110",
 2971 => "10110110",
 2972 => "00011001",
 2973 => "10001110",
 2974 => "10111011",
 2975 => "00110110",
 2976 => "00110111",
 2977 => "11100010",
 2978 => "00100001",
 2979 => "01100110",
 2980 => "11000000",
 2981 => "01010000",
 2982 => "00101101",
 2983 => "11010110",
 2984 => "01011001",
 2985 => "10001100",
 2986 => "10100100",
 2987 => "10101111",
 2988 => "01111010",
 2989 => "10001110",
 2990 => "11011111",
 2991 => "01000111",
 2992 => "01110001",
 2993 => "01101100",
 2994 => "10010001",
 2995 => "01010010",
 2996 => "11101010",
 2997 => "01101111",
 2998 => "11010011",
 2999 => "00110011",
 3000 => "10010111",
 3001 => "01110010",
 3002 => "11100101",
 3003 => "10001101",
 3004 => "11111000",
 3005 => "01101111",
 3006 => "10111000",
 3007 => "01000101",
 3008 => "10100110",
 3009 => "01011101",
 3010 => "00111111",
 3011 => "01111001",
 3012 => "10000100",
 3013 => "00011100",
 3014 => "10000100",
 3015 => "00110011",
 3016 => "00010010",
 3017 => "01000000",
 3018 => "11111010",
 3019 => "11010100",
 3020 => "10111101",
 3021 => "11011011",
 3022 => "11010000",
 3023 => "00111000",
 3024 => "10010011",
 3025 => "11001101",
 3026 => "01010111",
 3027 => "10001011",
 3028 => "10001000",
 3029 => "10000001",
 3030 => "01110110",
 3031 => "01000001",
 3032 => "11000101",
 3033 => "11001110",
 3034 => "00101101",
 3035 => "10111111",
 3036 => "01100011",
 3037 => "10100010",
 3038 => "01101001",
 3039 => "11010010",
 3040 => "00100110",
 3041 => "01010111",
 3042 => "01010100",
 3043 => "00101001",
 3044 => "11100011",
 3045 => "11011101",
 3046 => "00011000",
 3047 => "10001111",
 3048 => "11011111",
 3049 => "11111010",
 3050 => "01100111",
 3051 => "00001011",
 3052 => "01010111",
 3053 => "11011101",
 3054 => "10000101",
 3055 => "00111001",
 3056 => "11011100",
 3057 => "01100111",
 3058 => "01011000",
 3059 => "01011001",
 3060 => "11011111",
 3061 => "00001101",
 3062 => "00000101",
 3063 => "11010110",
 3064 => "11110111",
 3065 => "10110000",
 3066 => "00111111",
 3067 => "00111000",
 3068 => "11100111",
 3069 => "11101000",
 3070 => "01110100",
 3071 => "00101111",
 3072 => "11001101",
 3073 => "10110111",
 3074 => "01000111",
 3075 => "00001111",
 3076 => "00110110",
 3077 => "01100010",
 3078 => "11000010",
 3079 => "00011110",
 3080 => "10110000",
 3081 => "11100111",
 3082 => "10001100",
 3083 => "00001101",
 3084 => "00111010",
 3085 => "10000010",
 3086 => "00111111",
 3087 => "00010001",
 3088 => "00010111",
 3089 => "01110101",
 3090 => "10100010",
 3091 => "10111011",
 3092 => "00001100",
 3093 => "11111111",
 3094 => "10000111",
 3095 => "01111111",
 3096 => "01000001",
 3097 => "11111001",
 3098 => "11101100",
 3099 => "00010101",
 3100 => "01001111",
 3101 => "10000110",
 3102 => "10110101",
 3103 => "01100110",
 3104 => "11010001",
 3105 => "11001011",
 3106 => "00011000",
 3107 => "11110101",
 3108 => "10110111",
 3109 => "10111001",
 3110 => "01100101",
 3111 => "10011110",
 3112 => "01101001",
 3113 => "11000100",
 3114 => "01010100",
 3115 => "11100111",
 3116 => "00100010",
 3117 => "01000100",
 3118 => "01011100",
 3119 => "00000101",
 3120 => "01001101",
 3121 => "00010101",
 3122 => "11101111",
 3123 => "01100011",
 3124 => "11011011",
 3125 => "11100000",
 3126 => "10100011",
 3127 => "11000110",
 3128 => "10101010",
 3129 => "01111001",
 3130 => "01010101",
 3131 => "00100101",
 3132 => "11101101",
 3133 => "00000110",
 3134 => "11000110",
 3135 => "10001101",
 3136 => "00000100",
 3137 => "11111011",
 3138 => "00011111",
 3139 => "00000000",
 3140 => "00100000",
 3141 => "10010111",
 3142 => "11010011",
 3143 => "11111000",
 3144 => "01011010",
 3145 => "00011010",
 3146 => "11011100",
 3147 => "00010010",
 3148 => "10011001",
 3149 => "10111110",
 3150 => "01111110",
 3151 => "10001001",
 3152 => "11101110",
 3153 => "00110010",
 3154 => "10011011",
 3155 => "11011011",
 3156 => "11111010",
 3157 => "01110000",
 3158 => "11111111",
 3159 => "10111101",
 3160 => "00001011",
 3161 => "00000100",
 3162 => "11010001",
 3163 => "11001011",
 3164 => "00001110",
 3165 => "00010000",
 3166 => "01011101",
 3167 => "11000111",
 3168 => "11101100",
 3169 => "10010111",
 3170 => "01110001",
 3171 => "10010100",
 3172 => "11111000",
 3173 => "10000110",
 3174 => "00101000",
 3175 => "10001101",
 3176 => "00101010",
 3177 => "01110111",
 3178 => "00100110",
 3179 => "11010111",
 3180 => "00100011",
 3181 => "10000110",
 3182 => "00100100",
 3183 => "11000001",
 3184 => "10100111",
 3185 => "00000111",
 3186 => "01001010",
 3187 => "00101000",
 3188 => "00011111",
 3189 => "11000001",
 3190 => "00001001",
 3191 => "01111111",
 3192 => "01001110",
 3193 => "11010000",
 3194 => "11011010",
 3195 => "01110010",
 3196 => "01111111",
 3197 => "01000011",
 3198 => "10100001",
 3199 => "00011100",
 3200 => "11010000",
 3201 => "01001010",
 3202 => "11010011",
 3203 => "10101100",
 3204 => "10010111",
 3205 => "11010100",
 3206 => "11001111",
 3207 => "10100000",
 3208 => "01011110",
 3209 => "00011111",
 3210 => "01000101",
 3211 => "01011000",
 3212 => "10101011",
 3213 => "00010001",
 3214 => "10101101",
 3215 => "11110110",
 3216 => "00000110",
 3217 => "10111101",
 3218 => "01111101",
 3219 => "11111011",
 3220 => "00100000",
 3221 => "01000101",
 3222 => "00100111",
 3223 => "10100001",
 3224 => "00001111",
 3225 => "11100001",
 3226 => "10010100",
 3227 => "00100000",
 3228 => "11000101",
 3229 => "00100001",
 3230 => "10100001",
 3231 => "11011101",
 3232 => "10100101",
 3233 => "00011101",
 3234 => "11100001",
 3235 => "01000010",
 3236 => "10010010",
 3237 => "01010111",
 3238 => "10100011",
 3239 => "10011101",
 3240 => "10100010",
 3241 => "11101000",
 3242 => "11100011",
 3243 => "00011011",
 3244 => "00000001",
 3245 => "11100110",
 3246 => "01011010",
 3247 => "11110010",
 3248 => "10001110",
 3249 => "00100111",
 3250 => "11101011",
 3251 => "00000010",
 3252 => "11110110",
 3253 => "01001000",
 3254 => "01110111",
 3255 => "11001100",
 3256 => "10111110",
 3257 => "11101010",
 3258 => "10001001",
 3259 => "11101011",
 3260 => "10111110",
 3261 => "11011011",
 3262 => "10011111",
 3263 => "01000010",
 3264 => "10101111",
 3265 => "00111100",
 3266 => "10010111",
 3267 => "11110100",
 3268 => "11100000",
 3269 => "01110111",
 3270 => "00010100",
 3271 => "11010011",
 3272 => "01111001",
 3273 => "10000011",
 3274 => "10010111",
 3275 => "11100010",
 3276 => "10000110",
 3277 => "10000110",
 3278 => "10010000",
 3279 => "00111000",
 3280 => "01111010",
 3281 => "01110101",
 3282 => "01110101",
 3283 => "11111001",
 3284 => "00011101",
 3285 => "11110110",
 3286 => "00110000",
 3287 => "00001110",
 3288 => "11111011",
 3289 => "01101110",
 3290 => "00010101",
 3291 => "11110111",
 3292 => "01111010",
 3293 => "01100100",
 3294 => "11010001",
 3295 => "01110100",
 3296 => "00001001",
 3297 => "11000011",
 3298 => "00001111",
 3299 => "00010001",
 3300 => "01000011",
 3301 => "00110010",
 3302 => "00111110",
 3303 => "01101101",
 3304 => "00100100",
 3305 => "11000000",
 3306 => "00011010",
 3307 => "01000000",
 3308 => "10000111",
 3309 => "01011010",
 3310 => "00010101",
 3311 => "10010010",
 3312 => "11011010",
 3313 => "00111000",
 3314 => "01100111",
 3315 => "11111001",
 3316 => "11100010",
 3317 => "01110100",
 3318 => "10010000",
 3319 => "01100101",
 3320 => "00100010",
 3321 => "01011010",
 3322 => "10111101",
 3323 => "01000011",
 3324 => "11101001",
 3325 => "01011010",
 3326 => "00110100",
 3327 => "10001100",
 3328 => "00110001",
 3329 => "01011100",
 3330 => "00110000",
 3331 => "11100000",
 3332 => "10111000",
 3333 => "11000010",
 3334 => "00001100",
 3335 => "01111110",
 3336 => "10010001",
 3337 => "11000001",
 3338 => "01011001",
 3339 => "11000101",
 3340 => "10100111",
 3341 => "00011101",
 3342 => "10010010",
 3343 => "00010111",
 3344 => "01110001",
 3345 => "10010110",
 3346 => "00000100",
 3347 => "11110010",
 3348 => "01100010",
 3349 => "00000101",
 3350 => "10000011",
 3351 => "10011000",
 3352 => "01011000",
 3353 => "10101010",
 3354 => "01101110",
 3355 => "10100001",
 3356 => "11001000",
 3357 => "11011110",
 3358 => "10001101",
 3359 => "10001010",
 3360 => "11011101",
 3361 => "00011000",
 3362 => "10001101",
 3363 => "01100110",
 3364 => "01110100",
 3365 => "00110000",
 3366 => "11110010",
 3367 => "10111001",
 3368 => "11101010",
 3369 => "10100110",
 3370 => "10001001",
 3371 => "10001100",
 3372 => "01101011",
 3373 => "11100011",
 3374 => "00110100",
 3375 => "01000001",
 3376 => "10101101",
 3377 => "10011111",
 3378 => "01110011",
 3379 => "00100000",
 3380 => "11001100",
 3381 => "00111110",
 3382 => "11001110",
 3383 => "11100110",
 3384 => "10000100",
 3385 => "00001101",
 3386 => "00101011",
 3387 => "10011000",
 3388 => "10101010",
 3389 => "11111111",
 3390 => "11000010",
 3391 => "11100100",
 3392 => "00011000",
 3393 => "11101000",
 3394 => "00000001",
 3395 => "10110111",
 3396 => "00010010",
 3397 => "00101001",
 3398 => "11100110",
 3399 => "10010010",
 3400 => "01001010",
 3401 => "11000001",
 3402 => "00001011",
 3403 => "00011101",
 3404 => "10100011",
 3405 => "10100000",
 3406 => "00011110",
 3407 => "11100011",
 3408 => "11010011",
 3409 => "11010010",
 3410 => "01101110",
 3411 => "00011101",
 3412 => "11110100",
 3413 => "10000010",
 3414 => "00100010",
 3415 => "11010111",
 3416 => "10010100",
 3417 => "00001100",
 3418 => "11110110",
 3419 => "11011001",
 3420 => "01001000",
 3421 => "00000010",
 3422 => "00110111",
 3423 => "01111010",
 3424 => "10100001",
 3425 => "00111011",
 3426 => "11010011",
 3427 => "10110111",
 3428 => "11111100",
 3429 => "01101000",
 3430 => "00111100",
 3431 => "00011110",
 3432 => "01010011",
 3433 => "10111101",
 3434 => "01010011",
 3435 => "00110111",
 3436 => "11100100",
 3437 => "00101101",
 3438 => "11011101",
 3439 => "10000001",
 3440 => "10101010",
 3441 => "11010010",
 3442 => "01101010",
 3443 => "00011011",
 3444 => "00110000",
 3445 => "01011100",
 3446 => "11000010",
 3447 => "10110010",
 3448 => "11001010",
 3449 => "01111110",
 3450 => "11110011",
 3451 => "10000011",
 3452 => "10010001",
 3453 => "01010100",
 3454 => "00000111",
 3455 => "10011010",
 3456 => "11001101",
 3457 => "10011000",
 3458 => "10000111",
 3459 => "00101010",
 3460 => "00011101",
 3461 => "10110001",
 3462 => "11100001",
 3463 => "10100100",
 3464 => "00100011",
 3465 => "00000101",
 3466 => "01011100",
 3467 => "00010001",
 3468 => "11010000",
 3469 => "10110000",
 3470 => "01010101",
 3471 => "11101110",
 3472 => "11110110",
 3473 => "00110100",
 3474 => "00011001",
 3475 => "10100011",
 3476 => "10001011",
 3477 => "00111110",
 3478 => "11100111",
 3479 => "11110010",
 3480 => "10001000",
 3481 => "01010101",
 3482 => "01110101",
 3483 => "11010010",
 3484 => "11111011",
 3485 => "01100011",
 3486 => "00111111",
 3487 => "10001010",
 3488 => "00101100",
 3489 => "01100100",
 3490 => "10000100",
 3491 => "01000010",
 3492 => "00010110",
 3493 => "11000101",
 3494 => "11110111",
 3495 => "11110000",
 3496 => "00100011",
 3497 => "00101001",
 3498 => "01110100",
 3499 => "10011000",
 3500 => "00011010",
 3501 => "10110100",
 3502 => "00101001",
 3503 => "00101100",
 3504 => "10010010",
 3505 => "11010111",
 3506 => "11010111",
 3507 => "00100010",
 3508 => "01011010",
 3509 => "11111010",
 3510 => "11111111",
 3511 => "10110010",
 3512 => "10110010",
 3513 => "10000110",
 3514 => "10000000",
 3515 => "10111000",
 3516 => "00010011",
 3517 => "10001001",
 3518 => "10000001",
 3519 => "10101000",
 3520 => "00000101",
 3521 => "01010111",
 3522 => "11010011",
 3523 => "10111100",
 3524 => "10101010",
 3525 => "00100111",
 3526 => "11100111",
 3527 => "01000011",
 3528 => "11011101",
 3529 => "10110101",
 3530 => "01101001",
 3531 => "00100010",
 3532 => "10111001",
 3533 => "00011000",
 3534 => "11011111",
 3535 => "11011110",
 3536 => "11000110",
 3537 => "10100100",
 3538 => "10001111",
 3539 => "00100101",
 3540 => "11011011",
 3541 => "10101101",
 3542 => "00110001",
 3543 => "11001010",
 3544 => "10000110",
 3545 => "10101000",
 3546 => "00001111",
 3547 => "01101001",
 3548 => "10011011",
 3549 => "00111000",
 3550 => "11011111",
 3551 => "10101000",
 3552 => "11001101",
 3553 => "01011101",
 3554 => "00110000",
 3555 => "10010111",
 3556 => "01111101",
 3557 => "11001000",
 3558 => "11001111",
 3559 => "00101000",
 3560 => "10101010",
 3561 => "01110100",
 3562 => "00001110",
 3563 => "11001101",
 3564 => "01111101",
 3565 => "10100001",
 3566 => "11010111",
 3567 => "10110100",
 3568 => "00100111",
 3569 => "00010101",
 3570 => "01100011",
 3571 => "00111100",
 3572 => "01000010",
 3573 => "10111100",
 3574 => "01101010",
 3575 => "11001100",
 3576 => "01100010",
 3577 => "11101011",
 3578 => "11100101",
 3579 => "10000100",
 3580 => "10111011",
 3581 => "00011111",
 3582 => "10001001",
 3583 => "11111101",
 3584 => "10100110",
 3585 => "00111101",
 3586 => "01011010",
 3587 => "00111010",
 3588 => "11000001",
 3589 => "01011101",
 3590 => "11000110",
 3591 => "11010001",
 3592 => "10100000",
 3593 => "10110010",
 3594 => "11110100",
 3595 => "11101010",
 3596 => "10000000",
 3597 => "10100110",
 3598 => "10101001",
 3599 => "11100001",
 3600 => "01011101",
 3601 => "10111100",
 3602 => "01111010",
 3603 => "00001000",
 3604 => "11001101",
 3605 => "01110011",
 3606 => "00001100",
 3607 => "11010111",
 3608 => "11001001",
 3609 => "11001100",
 3610 => "11000110",
 3611 => "10000010",
 3612 => "00001001",
 3613 => "11111001",
 3614 => "00001011",
 3615 => "00110011",
 3616 => "01111011",
 3617 => "11101010",
 3618 => "10110101",
 3619 => "10111111",
 3620 => "00111111",
 3621 => "10001011",
 3622 => "11011011",
 3623 => "10011111",
 3624 => "11010101",
 3625 => "00000001",
 3626 => "11010011",
 3627 => "01101101",
 3628 => "00101001",
 3629 => "00111000",
 3630 => "01110000",
 3631 => "00101001",
 3632 => "11110110",
 3633 => "01010110",
 3634 => "01100001",
 3635 => "01100001",
 3636 => "00101111",
 3637 => "00010100",
 3638 => "11000110",
 3639 => "11011001",
 3640 => "10111110",
 3641 => "01110000",
 3642 => "01010001",
 3643 => "00000000",
 3644 => "11110011",
 3645 => "01110100",
 3646 => "11110011",
 3647 => "10011110",
 3648 => "11010000",
 3649 => "01000000",
 3650 => "01100110",
 3651 => "00100101",
 3652 => "10010101",
 3653 => "11101001",
 3654 => "11111001",
 3655 => "11100101",
 3656 => "00100011",
 3657 => "00010010",
 3658 => "10010101",
 3659 => "10010110",
 3660 => "01100100",
 3661 => "00001111",
 3662 => "01100000",
 3663 => "11010111",
 3664 => "01111111",
 3665 => "00000101",
 3666 => "00010100",
 3667 => "11011111",
 3668 => "10100001",
 3669 => "00100001",
 3670 => "01101111",
 3671 => "10100110",
 3672 => "00100101",
 3673 => "01011100",
 3674 => "11000000",
 3675 => "01010001",
 3676 => "10101111",
 3677 => "10110100",
 3678 => "10011101",
 3679 => "00000011",
 3680 => "11001000",
 3681 => "11100000",
 3682 => "10011011",
 3683 => "11010010",
 3684 => "01010011",
 3685 => "01110100",
 3686 => "11000110",
 3687 => "11010100",
 3688 => "10010101",
 3689 => "10000101",
 3690 => "01000010",
 3691 => "10000011",
 3692 => "01011000",
 3693 => "10111110",
 3694 => "11100011",
 3695 => "11011010",
 3696 => "01001011",
 3697 => "11111101",
 3698 => "11111001",
 3699 => "11011000",
 3700 => "01000110",
 3701 => "00001010",
 3702 => "00001111",
 3703 => "00000011",
 3704 => "00011011",
 3705 => "11100010",
 3706 => "11110001",
 3707 => "10011110",
 3708 => "10001101",
 3709 => "01110000",
 3710 => "00010111",
 3711 => "01011010",
 3712 => "11000011",
 3713 => "10100100",
 3714 => "10000110",
 3715 => "00101110",
 3716 => "00001001",
 3717 => "01000010",
 3718 => "10100010",
 3719 => "01100000",
 3720 => "01111111",
 3721 => "01000101",
 3722 => "00000000",
 3723 => "10100011",
 3724 => "11000001",
 3725 => "01001000",
 3726 => "11001010",
 3727 => "01100011",
 3728 => "00001101",
 3729 => "01101111",
 3730 => "00101001",
 3731 => "11001011",
 3732 => "01001011",
 3733 => "00110000",
 3734 => "01110001",
 3735 => "00000111",
 3736 => "10100111",
 3737 => "01001100",
 3738 => "01111011",
 3739 => "11100100",
 3740 => "00111001",
 3741 => "01000100",
 3742 => "00011110",
 3743 => "11110101",
 3744 => "10000000",
 3745 => "10101111",
 3746 => "00111111",
 3747 => "10011011",
 3748 => "01011110",
 3749 => "00000011",
 3750 => "11000101",
 3751 => "01011101",
 3752 => "10000000",
 3753 => "10111110",
 3754 => "00010110",
 3755 => "10111100",
 3756 => "10111001",
 3757 => "11101011",
 3758 => "00010100",
 3759 => "11011100",
 3760 => "01111100",
 3761 => "00011000",
 3762 => "00101100",
 3763 => "11011100",
 3764 => "11111001",
 3765 => "01111111",
 3766 => "10110011",
 3767 => "01110010",
 3768 => "10001101",
 3769 => "10001011",
 3770 => "01010010",
 3771 => "10001010",
 3772 => "00101100",
 3773 => "10100000",
 3774 => "01111111",
 3775 => "11110111",
 3776 => "01100000",
 3777 => "11001001",
 3778 => "10011010",
 3779 => "11001000",
 3780 => "00000010",
 3781 => "10111101",
 3782 => "10111000",
 3783 => "00010001",
 3784 => "00001101",
 3785 => "10110100",
 3786 => "00111111",
 3787 => "11010111",
 3788 => "00100101",
 3789 => "00010110",
 3790 => "01011101",
 3791 => "10000010",
 3792 => "10011110",
 3793 => "00111111",
 3794 => "00110111",
 3795 => "00011101",
 3796 => "10001111",
 3797 => "10001100",
 3798 => "11101100",
 3799 => "00001010",
 3800 => "01010110",
 3801 => "10001011",
 3802 => "01101001",
 3803 => "10011000",
 3804 => "00010010",
 3805 => "01000100",
 3806 => "00100110",
 3807 => "11110011",
 3808 => "00110110",
 3809 => "01011000",
 3810 => "11011011",
 3811 => "10101101",
 3812 => "00000000",
 3813 => "11000001",
 3814 => "01010011",
 3815 => "11100110",
 3816 => "11110010",
 3817 => "10111111",
 3818 => "11110101",
 3819 => "10100010",
 3820 => "11111110",
 3821 => "11111011",
 3822 => "10111011",
 3823 => "11101101",
 3824 => "01101101",
 3825 => "01010001",
 3826 => "10000010",
 3827 => "11011001",
 3828 => "00001001",
 3829 => "11000111",
 3830 => "11111001",
 3831 => "11110001",
 3832 => "10100010",
 3833 => "00010010",
 3834 => "01010000",
 3835 => "01111110",
 3836 => "10010100",
 3837 => "00111110",
 3838 => "11101110",
 3839 => "10001100",
 3840 => "00010000",
 3841 => "10111000",
 3842 => "11110011",
 3843 => "01000011",
 3844 => "00001110",
 3845 => "10011100",
 3846 => "11110100",
 3847 => "11001101",
 3848 => "00100110",
 3849 => "01000101",
 3850 => "11000001",
 3851 => "00111001",
 3852 => "11001010",
 3853 => "01101101",
 3854 => "01010101",
 3855 => "11001001",
 3856 => "00001100",
 3857 => "11000011",
 3858 => "01100101",
 3859 => "11011000",
 3860 => "00001100",
 3861 => "11000010",
 3862 => "00011000",
 3863 => "11000001",
 3864 => "11000100",
 3865 => "10000100",
 3866 => "00001111",
 3867 => "01101111",
 3868 => "10000000",
 3869 => "10101111",
 3870 => "10010011",
 3871 => "00100101",
 3872 => "10001100",
 3873 => "00110100",
 3874 => "00111010",
 3875 => "11001111",
 3876 => "00001100",
 3877 => "11110011",
 3878 => "00101001",
 3879 => "00100001",
 3880 => "10010010",
 3881 => "11101000",
 3882 => "01010011",
 3883 => "10101101",
 3884 => "01101111",
 3885 => "01101001",
 3886 => "10001101",
 3887 => "11011000",
 3888 => "10101000",
 3889 => "00000001",
 3890 => "00001011",
 3891 => "00000110",
 3892 => "11101111",
 3893 => "10110001",
 3894 => "11001001",
 3895 => "01101110",
 3896 => "01100000",
 3897 => "01000010",
 3898 => "01001000",
 3899 => "00110101",
 3900 => "10011010",
 3901 => "00100101",
 3902 => "00001001",
 3903 => "00110111",
 3904 => "01111011",
 3905 => "01101000",
 3906 => "10000011",
 3907 => "01101111",
 3908 => "10011101",
 3909 => "01100101",
 3910 => "11111001",
 3911 => "11110011",
 3912 => "00110110",
 3913 => "11100110",
 3914 => "11011001",
 3915 => "00000001",
 3916 => "11011111",
 3917 => "01001010",
 3918 => "11101111",
 3919 => "01100010",
 3920 => "00000011",
 3921 => "00101010",
 3922 => "01010110",
 3923 => "10101001",
 3924 => "10101011",
 3925 => "01011110",
 3926 => "00011011",
 3927 => "10101100",
 3928 => "01100111",
 3929 => "00101100",
 3930 => "10111100",
 3931 => "01110011",
 3932 => "00000011",
 3933 => "11010001",
 3934 => "00001111",
 3935 => "00010101",
 3936 => "11111100",
 3937 => "11101101",
 3938 => "00100000",
 3939 => "01101100",
 3940 => "00110010",
 3941 => "01010111",
 3942 => "00001101",
 3943 => "01001100",
 3944 => "01101110",
 3945 => "10011111",
 3946 => "11100011",
 3947 => "11001101",
 3948 => "10100100",
 3949 => "10101101",
 3950 => "10110110",
 3951 => "01101001",
 3952 => "01001001",
 3953 => "11100001",
 3954 => "01100101",
 3955 => "11000001",
 3956 => "00001101",
 3957 => "10101100",
 3958 => "00010110",
 3959 => "01101101",
 3960 => "00001110",
 3961 => "11101110",
 3962 => "01101011",
 3963 => "10100101",
 3964 => "10000101",
 3965 => "00111011",
 3966 => "01111101",
 3967 => "11000101",
 3968 => "00110011",
 3969 => "10010001",
 3970 => "10011101",
 3971 => "11001010",
 3972 => "11011001",
 3973 => "00110100",
 3974 => "01100111",
 3975 => "10100011",
 3976 => "11110011",
 3977 => "11000011",
 3978 => "11111011",
 3979 => "01101111",
 3980 => "00111111",
 3981 => "11100010",
 3982 => "01110100",
 3983 => "01100011",
 3984 => "11010011",
 3985 => "10010100",
 3986 => "11010111",
 3987 => "01101111",
 3988 => "00000101",
 3989 => "11101010",
 3990 => "01011110",
 3991 => "00011100",
 3992 => "11001000",
 3993 => "01110101",
 3994 => "01111011",
 3995 => "00111110",
 3996 => "11010100",
 3997 => "11001101",
 3998 => "11101111",
 3999 => "00111000",
 4000 => "00000000",
 4001 => "10110001",
 4002 => "10111110",
 4003 => "10001011",
 4004 => "10111000",
 4005 => "00101000",
 4006 => "00111111",
 4007 => "11101010",
 4008 => "01000000",
 4009 => "00100011",
 4010 => "11110111",
 4011 => "10001101",
 4012 => "00000101",
 4013 => "00011011",
 4014 => "10101001",
 4015 => "10111011",
 4016 => "10110010",
 4017 => "01100111",
 4018 => "11000000",
 4019 => "11110111",
 4020 => "00100010",
 4021 => "01111100",
 4022 => "10110010",
 4023 => "11001000",
 4024 => "11111110",
 4025 => "00010101",
 4026 => "10101000",
 4027 => "10001110",
 4028 => "00000101",
 4029 => "01100110",
 4030 => "10000100",
 4031 => "10011000",
 4032 => "10001110",
 4033 => "10101111",
 4034 => "01111001",
 4035 => "01100001",
 4036 => "01011010",
 4037 => "10100100",
 4038 => "00011011",
 4039 => "11101001",
 4040 => "11110011",
 4041 => "00110000",
 4042 => "10101110",
 4043 => "11111110",
 4044 => "10101100",
 4045 => "01100101",
 4046 => "10100001",
 4047 => "01011000",
 4048 => "00110010",
 4049 => "01001110",
 4050 => "00101010",
 4051 => "00000101",
 4052 => "11000000",
 4053 => "00001011",
 4054 => "00010111",
 4055 => "00110001",
 4056 => "11101000",
 4057 => "11010100",
 4058 => "00010101",
 4059 => "10110111",
 4060 => "10000001",
 4061 => "10111111",
 4062 => "00010100",
 4063 => "01000110",
 4064 => "11100111",
 4065 => "11100111",
 4066 => "01001001",
 4067 => "01101010",
 4068 => "01110100",
 4069 => "00100001",
 4070 => "10011010",
 4071 => "10101111",
 4072 => "10110110",
 4073 => "00000110",
 4074 => "00000100",
 4075 => "11100100",
 4076 => "11100011",
 4077 => "00000011",
 4078 => "11001010",
 4079 => "01010010",
 4080 => "01010111",
 4081 => "10100110",
 4082 => "01110000",
 4083 => "11101010",
 4084 => "10001011",
 4085 => "10100001",
 4086 => "10001000",
 4087 => "10011011",
 4088 => "00100110",
 4089 => "01101100",
 4090 => "01111101",
 4091 => "10100111",
 4092 => "00101010",
 4093 => "10110010",
 4094 => "01111011",
 4095 => "10110110",
 4096 => "00101101",
 4097 => "10100111",
 4098 => "10001101",
 4099 => "00111111",
 4100 => "01110100",
 4101 => "01010111",
 4102 => "01110111",
 4103 => "01000000",
 4104 => "01000000",
 4105 => "10100110",
 4106 => "10001111",
 4107 => "00100101",
 4108 => "01001010",
 4109 => "01111100",
 4110 => "11111110",
 4111 => "11100101",
 4112 => "11101101",
 4113 => "01001010",
 4114 => "11100110",
 4115 => "11101000",
 4116 => "00100100",
 4117 => "00111101",
 4118 => "10000001",
 4119 => "01010111",
 4120 => "11101101",
 4121 => "00110100",
 4122 => "11011101",
 4123 => "10011111",
 4124 => "11100110",
 4125 => "01111100",
 4126 => "10001000",
 4127 => "10110101",
 4128 => "11101110",
 4129 => "00000011",
 4130 => "11000100",
 4131 => "00000001",
 4132 => "00001001",
 4133 => "01100100",
 4134 => "01100100",
 4135 => "00010001",
 4136 => "11001010",
 4137 => "01010101",
 4138 => "11110111",
 4139 => "11011100",
 4140 => "10110000",
 4141 => "01111011",
 4142 => "11010000",
 4143 => "01101011",
 4144 => "11011011",
 4145 => "10001111",
 4146 => "00111111",
 4147 => "00100011",
 4148 => "01000001",
 4149 => "00011010",
 4150 => "01111101",
 4151 => "01100000",
 4152 => "10010000",
 4153 => "01010011",
 4154 => "11100011",
 4155 => "10101000",
 4156 => "00110100",
 4157 => "11000110",
 4158 => "10111011",
 4159 => "00110011",
 4160 => "10000101",
 4161 => "10100101",
 4162 => "10111100",
 4163 => "11001001",
 4164 => "11101101",
 4165 => "00111001",
 4166 => "11010000",
 4167 => "00111001",
 4168 => "00101001",
 4169 => "11010100",
 4170 => "10010000",
 4171 => "00000110",
 4172 => "00001111",
 4173 => "10111110",
 4174 => "01111010",
 4175 => "10101010",
 4176 => "11010101",
 4177 => "11111000",
 4178 => "10101000",
 4179 => "00000001",
 4180 => "01000111",
 4181 => "11010010",
 4182 => "10001101",
 4183 => "01111110",
 4184 => "00110000",
 4185 => "10100010",
 4186 => "10001101",
 4187 => "11111110",
 4188 => "11110101",
 4189 => "10000011",
 4190 => "00010010",
 4191 => "10000110",
 4192 => "01110010",
 4193 => "10110000",
 4194 => "11101011",
 4195 => "10001001",
 4196 => "01011001",
 4197 => "10100101",
 4198 => "10100011",
 4199 => "10000100",
 4200 => "01101000",
 4201 => "11111101",
 4202 => "00101111",
 4203 => "00010000",
 4204 => "00001100",
 4205 => "01100011",
 4206 => "11100111",
 4207 => "10111000",
 4208 => "11001001",
 4209 => "10011100",
 4210 => "01100011",
 4211 => "01111011",
 4212 => "01011110",
 4213 => "11110011",
 4214 => "00101110",
 4215 => "10100100",
 4216 => "11010011",
 4217 => "00111110",
 4218 => "01111111",
 4219 => "10100011",
 4220 => "11100111",
 4221 => "01101010",
 4222 => "10101001",
 4223 => "10110001",
 4224 => "10000100",
 4225 => "11110001",
 4226 => "11010110",
 4227 => "00001100",
 4228 => "10100100",
 4229 => "10011000",
 4230 => "00101001",
 4231 => "10001001",
 4232 => "10000111",
 4233 => "01111101",
 4234 => "00100101",
 4235 => "00110011",
 4236 => "00001100",
 4237 => "01001000",
 4238 => "11101100",
 4239 => "11111000",
 4240 => "00100100",
 4241 => "00011100",
 4242 => "01011001",
 4243 => "00101101",
 4244 => "10100011",
 4245 => "01101010",
 4246 => "11011111",
 4247 => "10111100",
 4248 => "11101111",
 4249 => "10111001",
 4250 => "01110000",
 4251 => "00010111",
 4252 => "11110011",
 4253 => "11111111",
 4254 => "01001011",
 4255 => "11100110",
 4256 => "11000001",
 4257 => "10101110",
 4258 => "00000111",
 4259 => "10010000",
 4260 => "10011110",
 4261 => "01000011",
 4262 => "10000001",
 4263 => "10011010",
 4264 => "10000011",
 4265 => "00000110",
 4266 => "11110101",
 4267 => "11100001",
 4268 => "00000001",
 4269 => "00010111",
 4270 => "00010011",
 4271 => "10101110",
 4272 => "10001111",
 4273 => "10111110",
 4274 => "11000101",
 4275 => "10111011",
 4276 => "10110111",
 4277 => "01101110",
 4278 => "11111110",
 4279 => "10001010",
 4280 => "10000000",
 4281 => "11011111",
 4282 => "01100110",
 4283 => "01111010",
 4284 => "11010110",
 4285 => "00110001",
 4286 => "00011111",
 4287 => "00101111",
 4288 => "00010011",
 4289 => "00010011",
 4290 => "11100100",
 4291 => "01010111",
 4292 => "10110011",
 4293 => "11101000",
 4294 => "11110100",
 4295 => "10110010",
 4296 => "01111010",
 4297 => "01100100",
 4298 => "11111101",
 4299 => "10111011",
 4300 => "00011111",
 4301 => "00010010",
 4302 => "01001110",
 4303 => "01110011",
 4304 => "01101000",
 4305 => "01100100",
 4306 => "11101010",
 4307 => "00010010",
 4308 => "11000010",
 4309 => "10011111",
 4310 => "10000000",
 4311 => "00100111",
 4312 => "11001111",
 4313 => "10011111",
 4314 => "00100110",
 4315 => "10100001",
 4316 => "01110000",
 4317 => "01010010",
 4318 => "11100001",
 4319 => "11100101",
 4320 => "11111100",
 4321 => "10011100",
 4322 => "11011110",
 4323 => "11110111",
 4324 => "00011110",
 4325 => "00110100",
 4326 => "11100110",
 4327 => "10100000",
 4328 => "10010010",
 4329 => "00110010",
 4330 => "00110101",
 4331 => "00001011",
 4332 => "11111001",
 4333 => "10101101",
 4334 => "10011000",
 4335 => "11010010",
 4336 => "01001110",
 4337 => "01000110",
 4338 => "10010001",
 4339 => "01111011",
 4340 => "00101110",
 4341 => "00011110",
 4342 => "00011001",
 4343 => "00000111",
 4344 => "00101100",
 4345 => "01000000",
 4346 => "11101011",
 4347 => "01111000",
 4348 => "00110001",
 4349 => "00010111",
 4350 => "00110001",
 4351 => "01001010",
 4352 => "00100100",
 4353 => "00001000",
 4354 => "01110111",
 4355 => "11000101",
 4356 => "01101000",
 4357 => "10000001",
 4358 => "00000111",
 4359 => "11100101",
 4360 => "01101100",
 4361 => "11001110",
 4362 => "11110110",
 4363 => "00000001",
 4364 => "01010100",
 4365 => "10000101",
 4366 => "00101111",
 4367 => "01100101",
 4368 => "10000100",
 4369 => "00111101",
 4370 => "10011001",
 4371 => "11000111",
 4372 => "00110000",
 4373 => "00110111",
 4374 => "11001001",
 4375 => "01010010",
 4376 => "10000001",
 4377 => "11100011",
 4378 => "01011111",
 4379 => "00111010",
 4380 => "11010010",
 4381 => "01100101",
 4382 => "01011110",
 4383 => "00101100",
 4384 => "11000101",
 4385 => "01000011",
 4386 => "10001001",
 4387 => "11011001",
 4388 => "01011101",
 4389 => "00010001",
 4390 => "00011110",
 4391 => "10001101",
 4392 => "11010111",
 4393 => "00000001",
 4394 => "10001010",
 4395 => "10110101",
 4396 => "10111111",
 4397 => "10110100",
 4398 => "00100110",
 4399 => "01100011",
 4400 => "00001101",
 4401 => "01101011",
 4402 => "11111110",
 4403 => "11011011",
 4404 => "11001101",
 4405 => "10001110",
 4406 => "00101111",
 4407 => "00010100",
 4408 => "10000011",
 4409 => "11000111",
 4410 => "01100010",
 4411 => "10011100",
 4412 => "10000001",
 4413 => "00101100",
 4414 => "10010101",
 4415 => "01110111",
 4416 => "00000000",
 4417 => "01111100",
 4418 => "10011000",
 4419 => "10000011",
 4420 => "00101001",
 4421 => "11001111",
 4422 => "00000100",
 4423 => "00001001",
 4424 => "00000101",
 4425 => "11011100",
 4426 => "00101010",
 4427 => "01000101",
 4428 => "01011110",
 4429 => "10111010",
 4430 => "10110101",
 4431 => "10100001",
 4432 => "10010111",
 4433 => "10011010",
 4434 => "01110010",
 4435 => "00111110",
 4436 => "10100001",
 4437 => "11101101",
 4438 => "01000101",
 4439 => "11011100",
 4440 => "00110011",
 4441 => "01011010",
 4442 => "11100111",
 4443 => "10011010",
 4444 => "11100000",
 4445 => "00100100",
 4446 => "11100101",
 4447 => "00000010",
 4448 => "01101000",
 4449 => "01110011",
 4450 => "11100010",
 4451 => "11010101",
 4452 => "10001010",
 4453 => "10000011",
 4454 => "11010110",
 4455 => "01111100",
 4456 => "11001100",
 4457 => "10100100",
 4458 => "01100100",
 4459 => "00010110",
 4460 => "10010001",
 4461 => "00010000",
 4462 => "01111101",
 4463 => "10110101",
 4464 => "01001100",
 4465 => "01001000",
 4466 => "11001101",
 4467 => "10111101",
 4468 => "10001011",
 4469 => "11110110",
 4470 => "01001111",
 4471 => "10101011",
 4472 => "01110111",
 4473 => "11000010",
 4474 => "10001111",
 4475 => "10110000",
 4476 => "10100100",
 4477 => "10111110",
 4478 => "10001010",
 4479 => "11110110",
 4480 => "01101110",
 4481 => "11100011",
 4482 => "11111000",
 4483 => "00111101",
 4484 => "01001000",
 4485 => "00000110",
 4486 => "10100101",
 4487 => "11110001",
 4488 => "10011110",
 4489 => "01100000",
 4490 => "00100010",
 4491 => "01101110",
 4492 => "10001111",
 4493 => "11111100",
 4494 => "11101001",
 4495 => "01000101",
 4496 => "00101011",
 4497 => "01001101",
 4498 => "10111001",
 4499 => "01000111",
 4500 => "10000100",
 4501 => "00000011",
 4502 => "10101111",
 4503 => "00000011",
 4504 => "10000000",
 4505 => "11101111",
 4506 => "00101100",
 4507 => "11101101",
 4508 => "10011010",
 4509 => "10000010",
 4510 => "10100111",
 4511 => "10010101",
 4512 => "11001010",
 4513 => "11111001",
 4514 => "10001001",
 4515 => "01110010",
 4516 => "10110011",
 4517 => "01001000",
 4518 => "11111101",
 4519 => "00011111",
 4520 => "01101011",
 4521 => "01110101",
 4522 => "11100111",
 4523 => "01101010",
 4524 => "11001111",
 4525 => "00000000",
 4526 => "01000010",
 4527 => "00011101",
 4528 => "00111101",
 4529 => "00100111",
 4530 => "10000011",
 4531 => "01111001",
 4532 => "10000001",
 4533 => "00000001",
 4534 => "10000000",
 4535 => "11110101",
 4536 => "00101001",
 4537 => "01000010",
 4538 => "10101110",
 4539 => "01111010",
 4540 => "01101011",
 4541 => "10101111",
 4542 => "01010110",
 4543 => "10001000",
 4544 => "00110000",
 4545 => "01001011",
 4546 => "10001101",
 4547 => "01111101",
 4548 => "11010100",
 4549 => "10000110",
 4550 => "10101001",
 4551 => "01110100",
 4552 => "11100111",
 4553 => "01010100",
 4554 => "01010111",
 4555 => "00001111",
 4556 => "11010101",
 4557 => "00110110",
 4558 => "00001011",
 4559 => "00101101",
 4560 => "11000100",
 4561 => "01000110",
 4562 => "11001011",
 4563 => "01000000",
 4564 => "10001011",
 4565 => "10001111",
 4566 => "10100110",
 4567 => "00011010",
 4568 => "01011000",
 4569 => "00110100",
 4570 => "01110011",
 4571 => "01000010",
 4572 => "00010010",
 4573 => "00011111",
 4574 => "00111010",
 4575 => "10110000",
 4576 => "00010101",
 4577 => "01110110",
 4578 => "11010110",
 4579 => "00110110",
 4580 => "11110011",
 4581 => "11011110",
 4582 => "11010101",
 4583 => "11001111",
 4584 => "11100111",
 4585 => "11110101",
 4586 => "11000011",
 4587 => "00111110",
 4588 => "01001101",
 4589 => "11000001",
 4590 => "10000001",
 4591 => "00101001",
 4592 => "11101101",
 4593 => "11011000",
 4594 => "00101010",
 4595 => "10000110",
 4596 => "01101011",
 4597 => "01111100",
 4598 => "01100001",
 4599 => "10110111",
 4600 => "01001011",
 4601 => "11001111",
 4602 => "01001001",
 4603 => "10011101",
 4604 => "01001110",
 4605 => "11100011",
 4606 => "11101100",
 4607 => "11100011",
 4608 => "00010100",
 4609 => "10010111",
 4610 => "01111011",
 4611 => "10101110",
 4612 => "11011110",
 4613 => "01111110",
 4614 => "00111001",
 4615 => "01000101",
 4616 => "10011000",
 4617 => "01111100",
 4618 => "11010001",
 4619 => "00011000",
 4620 => "01001010",
 4621 => "10110001",
 4622 => "11000001",
 4623 => "00010000",
 4624 => "00110010",
 4625 => "00111010",
 4626 => "10110101",
 4627 => "11000001",
 4628 => "01101000",
 4629 => "00010111",
 4630 => "01101000",
 4631 => "10010001",
 4632 => "11100010",
 4633 => "01010100",
 4634 => "10011101",
 4635 => "10010000",
 4636 => "11000100",
 4637 => "11000000",
 4638 => "11100011",
 4639 => "11100001",
 4640 => "11110010",
 4641 => "11110100",
 4642 => "10111000",
 4643 => "11011110",
 4644 => "11001101",
 4645 => "01000011",
 4646 => "00000111",
 4647 => "10111011",
 4648 => "10111110",
 4649 => "01100001",
 4650 => "00111100",
 4651 => "10001000",
 4652 => "10111110",
 4653 => "11100010",
 4654 => "10110000",
 4655 => "01011110",
 4656 => "11100000",
 4657 => "10100001",
 4658 => "10011101",
 4659 => "11010001",
 4660 => "01000011",
 4661 => "00011000",
 4662 => "10011101",
 4663 => "01110111",
 4664 => "00011011",
 4665 => "01100100",
 4666 => "10111000",
 4667 => "11110110",
 4668 => "11101101",
 4669 => "10101001",
 4670 => "00110000",
 4671 => "01101100",
 4672 => "01011010",
 4673 => "01100100",
 4674 => "01111010",
 4675 => "11010111",
 4676 => "00101000",
 4677 => "00110011",
 4678 => "00110101",
 4679 => "01100111",
 4680 => "10000010",
 4681 => "11001000",
 4682 => "10000011",
 4683 => "00110001",
 4684 => "00110000",
 4685 => "01101010",
 4686 => "00111110",
 4687 => "11110111",
 4688 => "01001010",
 4689 => "11110001",
 4690 => "11001100",
 4691 => "10000001",
 4692 => "00101001",
 4693 => "11111000",
 4694 => "10110100",
 4695 => "00001110",
 4696 => "01110101",
 4697 => "00001000",
 4698 => "10001000",
 4699 => "01110100",
 4700 => "00000000",
 4701 => "00000000",
 4702 => "00011001",
 4703 => "00111110",
 4704 => "11001010",
 4705 => "11110110",
 4706 => "10111101",
 4707 => "10001011",
 4708 => "11011110",
 4709 => "01001001",
 4710 => "11011000",
 4711 => "00111010",
 4712 => "10001101",
 4713 => "00101111",
 4714 => "10101111",
 4715 => "11110000",
 4716 => "11010010",
 4717 => "00011010",
 4718 => "01100000",
 4719 => "11000100",
 4720 => "11000001",
 4721 => "01010101",
 4722 => "00010000",
 4723 => "10001000",
 4724 => "01001000",
 4725 => "01101100",
 4726 => "11100111",
 4727 => "10010100",
 4728 => "01111010",
 4729 => "00101101",
 4730 => "00010110",
 4731 => "11010100",
 4732 => "10000001",
 4733 => "10010011",
 4734 => "00100111",
 4735 => "10011011",
 4736 => "10010011",
 4737 => "01010111",
 4738 => "01110001",
 4739 => "01011010",
 4740 => "00001011",
 4741 => "11111011",
 4742 => "00011000",
 4743 => "01010011",
 4744 => "10100010",
 4745 => "11110010",
 4746 => "01000011",
 4747 => "10010111",
 4748 => "00011110",
 4749 => "10001000",
 4750 => "00100001",
 4751 => "00101011",
 4752 => "00011111",
 4753 => "00011110",
 4754 => "01001011",
 4755 => "01010010",
 4756 => "01011011",
 4757 => "01101001",
 4758 => "11000011",
 4759 => "01100011",
 4760 => "00101101",
 4761 => "01001010",
 4762 => "11111000",
 4763 => "01010000",
 4764 => "10000101",
 4765 => "11101010",
 4766 => "11000110",
 4767 => "01111100",
 4768 => "01111011",
 4769 => "10001001",
 4770 => "11001110",
 4771 => "00011010",
 4772 => "01000110",
 4773 => "11111011",
 4774 => "00101010",
 4775 => "00010111",
 4776 => "00111101",
 4777 => "11000110",
 4778 => "01001001",
 4779 => "11010101",
 4780 => "01110001",
 4781 => "01010001",
 4782 => "01111101",
 4783 => "11001011",
 4784 => "01110001",
 4785 => "01100001",
 4786 => "00011001",
 4787 => "01100010",
 4788 => "00101001",
 4789 => "11100010",
 4790 => "01100111",
 4791 => "00000011",
 4792 => "10111001",
 4793 => "10101100",
 4794 => "00111010",
 4795 => "01100000",
 4796 => "10001010",
 4797 => "01100011",
 4798 => "10010100",
 4799 => "11110000",
 4800 => "10011111",
 4801 => "01101100",
 4802 => "11001111",
 4803 => "01000000",
 4804 => "01010100",
 4805 => "00100101",
 4806 => "11001010",
 4807 => "11000100",
 4808 => "11011011",
 4809 => "10100010",
 4810 => "10011010",
 4811 => "10011100",
 4812 => "10000001",
 4813 => "10011101",
 4814 => "11010111",
 4815 => "11001111",
 4816 => "00010001",
 4817 => "11011000",
 4818 => "11011100",
 4819 => "00100001",
 4820 => "01101101",
 4821 => "00111111",
 4822 => "10011111",
 4823 => "01110101",
 4824 => "11010001",
 4825 => "00001000",
 4826 => "00000111",
 4827 => "10010000",
 4828 => "00101010",
 4829 => "11000011",
 4830 => "11001000",
 4831 => "01100011",
 4832 => "11011111",
 4833 => "11010010",
 4834 => "01000101",
 4835 => "00111000",
 4836 => "10010000",
 4837 => "01011100",
 4838 => "00100000",
 4839 => "11101100",
 4840 => "11100111",
 4841 => "10101110",
 4842 => "01010010",
 4843 => "01100100",
 4844 => "11110100",
 4845 => "01101100",
 4846 => "01101110",
 4847 => "11100110",
 4848 => "00010101",
 4849 => "11000010",
 4850 => "10001101",
 4851 => "01101001",
 4852 => "01010010",
 4853 => "00110001",
 4854 => "11000111",
 4855 => "10011010",
 4856 => "10101000",
 4857 => "00011101",
 4858 => "10100011",
 4859 => "10111111",
 4860 => "10000111",
 4861 => "00111101",
 4862 => "00111101",
 4863 => "11101100",
 4864 => "11000101",
 4865 => "10000001",
 4866 => "01010111",
 4867 => "10011100",
 4868 => "11101010",
 4869 => "11000001",
 4870 => "01011111",
 4871 => "10101000",
 4872 => "11111100",
 4873 => "01011110",
 4874 => "00111011",
 4875 => "10100110",
 4876 => "01010001",
 4877 => "00110001",
 4878 => "01000000",
 4879 => "10100010",
 4880 => "10010011",
 4881 => "01011100",
 4882 => "10111100",
 4883 => "01011101",
 4884 => "10010111",
 4885 => "11101110",
 4886 => "10100110",
 4887 => "11111001",
 4888 => "00000111",
 4889 => "00101101",
 4890 => "10101010",
 4891 => "01001010",
 4892 => "00110100",
 4893 => "11101000",
 4894 => "11000100",
 4895 => "10111101",
 4896 => "11000011",
 4897 => "11110011",
 4898 => "11011010",
 4899 => "11101001",
 4900 => "01100101",
 4901 => "11010000",
 4902 => "00000111",
 4903 => "01010110",
 4904 => "11110111",
 4905 => "00010111",
 4906 => "00011101",
 4907 => "11001001",
 4908 => "11100011",
 4909 => "00001100",
 4910 => "11101100",
 4911 => "11011001",
 4912 => "11110110",
 4913 => "11001000",
 4914 => "11111111",
 4915 => "01110100",
 4916 => "11011000",
 4917 => "11100101",
 4918 => "01001001",
 4919 => "01001100",
 4920 => "11111111",
 4921 => "00111000",
 4922 => "10100001",
 4923 => "01111001",
 4924 => "00101010",
 4925 => "11011001",
 4926 => "00100011",
 4927 => "11011011",
 4928 => "11100110",
 4929 => "00110010",
 4930 => "11000001",
 4931 => "11000111",
 4932 => "11110100",
 4933 => "01000110",
 4934 => "11111010",
 4935 => "00000100",
 4936 => "10011100",
 4937 => "10011010",
 4938 => "01010100",
 4939 => "01111111",
 4940 => "00010110",
 4941 => "11010010",
 4942 => "10110111",
 4943 => "10010111",
 4944 => "00101110",
 4945 => "11011111",
 4946 => "11110111",
 4947 => "01100000",
 4948 => "01101011",
 4949 => "10011100",
 4950 => "11000111",
 4951 => "10000000",
 4952 => "11110101",
 4953 => "00100111",
 4954 => "11111001",
 4955 => "11111111",
 4956 => "00010011",
 4957 => "11000110",
 4958 => "11000101",
 4959 => "01110010",
 4960 => "10011011",
 4961 => "01000110",
 4962 => "11110100",
 4963 => "01011010",
 4964 => "10110001",
 4965 => "10100001",
 4966 => "11011001",
 4967 => "11110101",
 4968 => "11101110",
 4969 => "10101110",
 4970 => "10100111",
 4971 => "00101011",
 4972 => "10010101",
 4973 => "01011110",
 4974 => "10000000",
 4975 => "10011111",
 4976 => "10010011",
 4977 => "01001101",
 4978 => "10100000",
 4979 => "10100011",
 4980 => "10010111",
 4981 => "01001101",
 4982 => "11010101",
 4983 => "11110000",
 4984 => "00100101",
 4985 => "11000011",
 4986 => "00000101",
 4987 => "01000111",
 4988 => "10111100",
 4989 => "10100010",
 4990 => "11100111",
 4991 => "10111110",
 4992 => "00001000",
 4993 => "10100111",
 4994 => "10110000",
 4995 => "10010011",
 4996 => "11001011",
 4997 => "00111000",
 4998 => "11010100",
 4999 => "00111011",
 5000 => "11010111",
 5001 => "01101111",
 5002 => "00111001",
 5003 => "00110001",
 5004 => "11011100",
 5005 => "10110001",
 5006 => "01101111",
 5007 => "00001000",
 5008 => "01110001",
 5009 => "11101111",
 5010 => "11001100",
 5011 => "11010111",
 5012 => "11001101",
 5013 => "10000010",
 5014 => "00101000",
 5015 => "10111110",
 5016 => "10001110",
 5017 => "11011110",
 5018 => "11001111",
 5019 => "01010101",
 5020 => "00101101",
 5021 => "10001111",
 5022 => "10101100",
 5023 => "00010010",
 5024 => "00100111",
 5025 => "10100011",
 5026 => "11101001",
 5027 => "10010110",
 5028 => "10110000",
 5029 => "10100101",
 5030 => "00101000",
 5031 => "00101001",
 5032 => "01001101",
 5033 => "10010010",
 5034 => "11011111",
 5035 => "11111110",
 5036 => "00111100",
 5037 => "01001001",
 5038 => "11001010",
 5039 => "00101100",
 5040 => "00111100",
 5041 => "00001111",
 5042 => "01010010",
 5043 => "11111010",
 5044 => "10000110",
 5045 => "10011001",
 5046 => "10010001",
 5047 => "10100101",
 5048 => "10110010",
 5049 => "10011101",
 5050 => "10110001",
 5051 => "00000111",
 5052 => "00000010",
 5053 => "00111010",
 5054 => "01010110",
 5055 => "11110111",
 5056 => "01001000",
 5057 => "11101111",
 5058 => "10110001",
 5059 => "00101000",
 5060 => "00010101",
 5061 => "00000101",
 5062 => "11110110",
 5063 => "00111000",
 5064 => "11000000",
 5065 => "01111001",
 5066 => "00110011",
 5067 => "11101000",
 5068 => "00110110",
 5069 => "00111110",
 5070 => "10100001",
 5071 => "01001101",
 5072 => "01101111",
 5073 => "11111001",
 5074 => "11101011",
 5075 => "11110011",
 5076 => "00110101",
 5077 => "00010110",
 5078 => "11100111",
 5079 => "01100011",
 5080 => "00001111",
 5081 => "11111100",
 5082 => "00110010",
 5083 => "11011000",
 5084 => "01001011",
 5085 => "11010000",
 5086 => "01111000",
 5087 => "00000101",
 5088 => "01001101",
 5089 => "10100011",
 5090 => "10100011",
 5091 => "00101100",
 5092 => "01000001",
 5093 => "00010001",
 5094 => "00011001",
 5095 => "10111001",
 5096 => "00010001",
 5097 => "00010101",
 5098 => "11110011",
 5099 => "10101000",
 5100 => "10010110",
 5101 => "10101011",
 5102 => "10010110",
 5103 => "10101111",
 5104 => "11100100",
 5105 => "00010101",
 5106 => "01100110",
 5107 => "00111110",
 5108 => "10111011",
 5109 => "00011100",
 5110 => "11100110",
 5111 => "10010100",
 5112 => "11010110",
 5113 => "00101101",
 5114 => "01111111",
 5115 => "00001110",
 5116 => "10110100",
 5117 => "10011010",
 5118 => "00001110",
 5119 => "00010100",
 5120 => "00111011",
 5121 => "00110111",
 5122 => "10001111",
 5123 => "10111101",
 5124 => "01100100",
 5125 => "11010111",
 5126 => "01010101",
 5127 => "10000100",
 5128 => "11110100",
 5129 => "01011110",
 5130 => "10010100",
 5131 => "01111001",
 5132 => "11100001",
 5133 => "00101110",
 5134 => "00110001",
 5135 => "00000001",
 5136 => "00011010",
 5137 => "00100010",
 5138 => "10100111",
 5139 => "00101100",
 5140 => "11011000",
 5141 => "10001101",
 5142 => "00100111",
 5143 => "10110111",
 5144 => "10111101",
 5145 => "11100110",
 5146 => "10110001",
 5147 => "10110010",
 5148 => "11000010",
 5149 => "01111001",
 5150 => "11000011",
 5151 => "01111100",
 5152 => "10110010",
 5153 => "00100110",
 5154 => "10111100",
 5155 => "01100000",
 5156 => "01001111",
 5157 => "11001101",
 5158 => "01011010",
 5159 => "10100101",
 5160 => "01001010",
 5161 => "00100010",
 5162 => "11001110",
 5163 => "11001001",
 5164 => "01011101",
 5165 => "11000100",
 5166 => "01100100",
 5167 => "00001111",
 5168 => "01000111",
 5169 => "11000001",
 5170 => "11101001",
 5171 => "11010000",
 5172 => "11011000",
 5173 => "00011010",
 5174 => "11010101",
 5175 => "11001001",
 5176 => "10011000",
 5177 => "00101010",
 5178 => "10000010",
 5179 => "11101101",
 5180 => "00010101",
 5181 => "01010100",
 5182 => "10100011",
 5183 => "01110101",
 5184 => "11110010",
 5185 => "11011001",
 5186 => "11001000",
 5187 => "10010000",
 5188 => "01111100",
 5189 => "00110101",
 5190 => "01011000",
 5191 => "01100011",
 5192 => "00111110",
 5193 => "10010101",
 5194 => "01111000",
 5195 => "00101111",
 5196 => "10111010",
 5197 => "00010010",
 5198 => "01101001",
 5199 => "00010111",
 5200 => "11101100",
 5201 => "01010010",
 5202 => "11111001",
 5203 => "11101010",
 5204 => "11111010",
 5205 => "00101000",
 5206 => "01101100",
 5207 => "11001000",
 5208 => "00011100",
 5209 => "11010111",
 5210 => "11101011",
 5211 => "01000010",
 5212 => "11111110",
 5213 => "00000010",
 5214 => "00111101",
 5215 => "00110111",
 5216 => "10010001",
 5217 => "11011111",
 5218 => "00001110",
 5219 => "10010110",
 5220 => "00101000",
 5221 => "10000100",
 5222 => "10011111",
 5223 => "01111001",
 5224 => "00100010",
 5225 => "10101101",
 5226 => "00001100",
 5227 => "11001110",
 5228 => "11000001",
 5229 => "10000101",
 5230 => "11000101",
 5231 => "11011011",
 5232 => "10101101",
 5233 => "01111011",
 5234 => "01010100",
 5235 => "00011110",
 5236 => "00000110",
 5237 => "01111001",
 5238 => "11101011",
 5239 => "01110011",
 5240 => "01001001",
 5241 => "10101000",
 5242 => "00110111",
 5243 => "11000101",
 5244 => "11001111",
 5245 => "00111000",
 5246 => "00010010",
 5247 => "01010100",
 5248 => "01111111",
 5249 => "11111011",
 5250 => "11110110",
 5251 => "11010010",
 5252 => "10001000",
 5253 => "11001001",
 5254 => "11111001",
 5255 => "00000101",
 5256 => "11110001",
 5257 => "01011100",
 5258 => "01101100",
 5259 => "00101100",
 5260 => "00010110",
 5261 => "11101000",
 5262 => "10110110",
 5263 => "00000001",
 5264 => "10100100",
 5265 => "11110110",
 5266 => "11000000",
 5267 => "10100100",
 5268 => "11100101",
 5269 => "11101110",
 5270 => "10111000",
 5271 => "11001101",
 5272 => "00010001",
 5273 => "10110101",
 5274 => "01110001",
 5275 => "00100101",
 5276 => "01110110",
 5277 => "10111001",
 5278 => "10011101",
 5279 => "01101111",
 5280 => "11000011",
 5281 => "11100101",
 5282 => "00001010",
 5283 => "01000101",
 5284 => "01001000",
 5285 => "10001000",
 5286 => "11110110",
 5287 => "10111101",
 5288 => "11001101",
 5289 => "10101110",
 5290 => "10001110",
 5291 => "01001111",
 5292 => "00011000",
 5293 => "10000010",
 5294 => "10010011",
 5295 => "11010011",
 5296 => "01101110",
 5297 => "10011111",
 5298 => "10000000",
 5299 => "10100100",
 5300 => "11110001",
 5301 => "00111011",
 5302 => "01011110",
 5303 => "11000110",
 5304 => "11010000",
 5305 => "10101111",
 5306 => "10010011",
 5307 => "01110011",
 5308 => "11101001",
 5309 => "01010110",
 5310 => "01010110",
 5311 => "10010000",
 5312 => "01010001",
 5313 => "11010000",
 5314 => "01000010",
 5315 => "11100001",
 5316 => "01001001",
 5317 => "11100001",
 5318 => "01011000",
 5319 => "11000101",
 5320 => "10011100",
 5321 => "01010110",
 5322 => "01011000",
 5323 => "01100111",
 5324 => "11110100",
 5325 => "11100000",
 5326 => "00010111",
 5327 => "11010110",
 5328 => "10110101",
 5329 => "10000101",
 5330 => "10000001",
 5331 => "01010100",
 5332 => "00001101",
 5333 => "11000001",
 5334 => "00011010",
 5335 => "01001101",
 5336 => "10111010",
 5337 => "01010110",
 5338 => "11001111",
 5339 => "00100111",
 5340 => "00010000",
 5341 => "00110011",
 5342 => "11110101",
 5343 => "10110010",
 5344 => "11011100",
 5345 => "11010101",
 5346 => "10111010",
 5347 => "00100110",
 5348 => "11011111",
 5349 => "00111110",
 5350 => "01110001",
 5351 => "11010011",
 5352 => "01011011",
 5353 => "11011101",
 5354 => "00011010",
 5355 => "10011011",
 5356 => "11000001",
 5357 => "01010110",
 5358 => "11011111",
 5359 => "00010001",
 5360 => "01111110",
 5361 => "01110010",
 5362 => "10011100",
 5363 => "00100100",
 5364 => "01110100",
 5365 => "10110101",
 5366 => "10011100",
 5367 => "01010111",
 5368 => "10010100",
 5369 => "01001100",
 5370 => "00101011",
 5371 => "10011010",
 5372 => "10001100",
 5373 => "10001001",
 5374 => "11001011",
 5375 => "00110111",
 5376 => "01010110",
 5377 => "11101110",
 5378 => "10101111",
 5379 => "11010110",
 5380 => "01010001",
 5381 => "11010100",
 5382 => "11111001",
 5383 => "01001100",
 5384 => "10100111",
 5385 => "01000000",
 5386 => "01011001",
 5387 => "01101101",
 5388 => "10101100",
 5389 => "01100011",
 5390 => "01010010",
 5391 => "01001001",
 5392 => "10101111",
 5393 => "10000000",
 5394 => "00101110",
 5395 => "00000110",
 5396 => "01101101",
 5397 => "11101101",
 5398 => "10011101",
 5399 => "11101010",
 5400 => "11100101",
 5401 => "10011110",
 5402 => "00110011",
 5403 => "11111000",
 5404 => "00010111",
 5405 => "01010101",
 5406 => "11010101",
 5407 => "01011111",
 5408 => "00010111",
 5409 => "11100101",
 5410 => "01010001",
 5411 => "01101001",
 5412 => "01111001",
 5413 => "11100111",
 5414 => "00100110",
 5415 => "01101011",
 5416 => "10001100",
 5417 => "01111111",
 5418 => "10100001",
 5419 => "10011110",
 5420 => "10011011",
 5421 => "10111110",
 5422 => "00001101",
 5423 => "00111111",
 5424 => "01000111",
 5425 => "01100000",
 5426 => "00000001",
 5427 => "01111000",
 5428 => "11100011",
 5429 => "01010101",
 5430 => "00000000",
 5431 => "10000110",
 5432 => "11101011",
 5433 => "00100101",
 5434 => "00011100",
 5435 => "10110011",
 5436 => "11100010",
 5437 => "00110111",
 5438 => "00101001",
 5439 => "01100000",
 5440 => "00011001",
 5441 => "11111000",
 5442 => "01101111",
 5443 => "01011000",
 5444 => "10011111",
 5445 => "10100001",
 5446 => "00101101",
 5447 => "00110110",
 5448 => "11101110",
 5449 => "01110101",
 5450 => "10110011",
 5451 => "00101101",
 5452 => "00110111",
 5453 => "00011000",
 5454 => "01100110",
 5455 => "10001110",
 5456 => "00010101",
 5457 => "01010010",
 5458 => "00000101",
 5459 => "10110001",
 5460 => "11111100",
 5461 => "10000001",
 5462 => "11110111",
 5463 => "11001010",
 5464 => "11010100",
 5465 => "01010100",
 5466 => "01011101",
 5467 => "10101111",
 5468 => "00110001",
 5469 => "11000101",
 5470 => "00110100",
 5471 => "11100001",
 5472 => "10100110",
 5473 => "01011011",
 5474 => "01111111",
 5475 => "00110110",
 5476 => "00100101",
 5477 => "01000000",
 5478 => "00100010",
 5479 => "01010001",
 5480 => "01001001",
 5481 => "10001010",
 5482 => "01101011",
 5483 => "11001011",
 5484 => "01000000",
 5485 => "01111101",
 5486 => "10111010",
 5487 => "00101011",
 5488 => "11100010",
 5489 => "11000001",
 5490 => "00110011",
 5491 => "01001110",
 5492 => "00001010",
 5493 => "00101000",
 5494 => "11110011",
 5495 => "01001111",
 5496 => "01101001",
 5497 => "00100010",
 5498 => "00110100",
 5499 => "00000100",
 5500 => "10111011",
 5501 => "11010111",
 5502 => "10101000",
 5503 => "00001011",
 5504 => "01001100",
 5505 => "01110000",
 5506 => "11101011",
 5507 => "10110010",
 5508 => "10010110",
 5509 => "00011111",
 5510 => "11011111",
 5511 => "00000101",
 5512 => "10011111",
 5513 => "01000111",
 5514 => "00110111",
 5515 => "00110111",
 5516 => "11111011",
 5517 => "01110010",
 5518 => "10000011",
 5519 => "11110000",
 5520 => "10000001",
 5521 => "11111101",
 5522 => "00101011",
 5523 => "11000011",
 5524 => "11010010",
 5525 => "01000001",
 5526 => "00101110",
 5527 => "00001010",
 5528 => "00001010",
 5529 => "10100010",
 5530 => "10111110",
 5531 => "11000010",
 5532 => "11010101",
 5533 => "11100001",
 5534 => "11010011",
 5535 => "00011111",
 5536 => "10000100",
 5537 => "00101111",
 5538 => "10111100",
 5539 => "10010001",
 5540 => "10110010",
 5541 => "00101100",
 5542 => "11000100",
 5543 => "10010111",
 5544 => "01111001",
 5545 => "10110010",
 5546 => "01000100",
 5547 => "00010110",
 5548 => "01000100",
 5549 => "01110010",
 5550 => "10010111",
 5551 => "00110000",
 5552 => "11010111",
 5553 => "11101111",
 5554 => "10100000",
 5555 => "10100010",
 5556 => "00011001",
 5557 => "10011000",
 5558 => "01110001",
 5559 => "10010100",
 5560 => "11001100",
 5561 => "01011101",
 5562 => "10101111",
 5563 => "01110000",
 5564 => "00001000",
 5565 => "10111001",
 5566 => "01000100",
 5567 => "11100110",
 5568 => "00011111",
 5569 => "10010000",
 5570 => "01010111",
 5571 => "10110001",
 5572 => "11111110",
 5573 => "10110000",
 5574 => "11011011",
 5575 => "11101111",
 5576 => "01000111",
 5577 => "01010000",
 5578 => "00010010",
 5579 => "11011010",
 5580 => "11110000",
 5581 => "11000011",
 5582 => "10010100",
 5583 => "00001101",
 5584 => "11000111",
 5585 => "11011100",
 5586 => "00001110",
 5587 => "01101000",
 5588 => "00100010",
 5589 => "11011000",
 5590 => "10010100",
 5591 => "10101000",
 5592 => "00110001",
 5593 => "10100101",
 5594 => "10010101",
 5595 => "01101110",
 5596 => "11111011",
 5597 => "10101001",
 5598 => "10110011",
 5599 => "10000001",
 5600 => "01011011",
 5601 => "00000100",
 5602 => "00110011",
 5603 => "11010001",
 5604 => "11110101",
 5605 => "11001111",
 5606 => "01010000",
 5607 => "01000001",
 5608 => "01101000",
 5609 => "11110111",
 5610 => "00010110",
 5611 => "11011110",
 5612 => "10111110",
 5613 => "01111101",
 5614 => "11100011",
 5615 => "00000110",
 5616 => "11001001",
 5617 => "10010011",
 5618 => "00111100",
 5619 => "01001011",
 5620 => "01101001",
 5621 => "00010110",
 5622 => "01011111",
 5623 => "10100010",
 5624 => "00000001",
 5625 => "10001001",
 5626 => "00101010",
 5627 => "11011001",
 5628 => "01111101",
 5629 => "00101100",
 5630 => "01111000",
 5631 => "00011111",
 5632 => "01001000",
 5633 => "00100011",
 5634 => "10000010",
 5635 => "11110111",
 5636 => "00101000",
 5637 => "10100001",
 5638 => "00110110",
 5639 => "10001000",
 5640 => "01001110",
 5641 => "01001000",
 5642 => "11011101",
 5643 => "10110111",
 5644 => "10110100",
 5645 => "01100000",
 5646 => "11100101",
 5647 => "00101111",
 5648 => "10110001",
 5649 => "01111000",
 5650 => "11100000",
 5651 => "01001000",
 5652 => "00100100",
 5653 => "01000011",
 5654 => "00000011",
 5655 => "00101101",
 5656 => "11101100",
 5657 => "10110010",
 5658 => "11111101",
 5659 => "01100011",
 5660 => "00010010",
 5661 => "01011011",
 5662 => "01001110",
 5663 => "00011101",
 5664 => "00000000",
 5665 => "11111110",
 5666 => "01110011",
 5667 => "01100001",
 5668 => "11011000",
 5669 => "11111100",
 5670 => "00001101",
 5671 => "11100010",
 5672 => "10111101",
 5673 => "11010111",
 5674 => "11100000",
 5675 => "00101000",
 5676 => "10010100",
 5677 => "11110101",
 5678 => "11011011",
 5679 => "01001011",
 5680 => "11001000",
 5681 => "11101000",
 5682 => "10110111",
 5683 => "01101110",
 5684 => "00001010",
 5685 => "11010000",
 5686 => "00100111",
 5687 => "10110101",
 5688 => "00000110",
 5689 => "01110111",
 5690 => "01000101",
 5691 => "01010100",
 5692 => "00111111",
 5693 => "01000000",
 5694 => "00110111",
 5695 => "10100111",
 5696 => "10101010",
 5697 => "00000010",
 5698 => "01100110",
 5699 => "10110111",
 5700 => "01101010",
 5701 => "01001110",
 5702 => "01001010",
 5703 => "10011000",
 5704 => "01111111",
 5705 => "01000001",
 5706 => "10000111",
 5707 => "00010111",
 5708 => "00001100",
 5709 => "00111010",
 5710 => "10110101",
 5711 => "01111111",
 5712 => "11010000",
 5713 => "10000000",
 5714 => "00010110",
 5715 => "00010110",
 5716 => "11010111",
 5717 => "01100001",
 5718 => "01001110",
 5719 => "11100011",
 5720 => "01001111",
 5721 => "10000101",
 5722 => "00101110",
 5723 => "10000000",
 5724 => "10011111",
 5725 => "01110001",
 5726 => "00111000",
 5727 => "00111110",
 5728 => "00110011",
 5729 => "00011011",
 5730 => "11001101",
 5731 => "11101000",
 5732 => "00101000",
 5733 => "00110111",
 5734 => "10100010",
 5735 => "01100011",
 5736 => "11101110",
 5737 => "10010010",
 5738 => "10111100",
 5739 => "01001011",
 5740 => "10111101",
 5741 => "01111000",
 5742 => "00101001",
 5743 => "11100100",
 5744 => "10100100",
 5745 => "11010001",
 5746 => "10111001",
 5747 => "00011000",
 5748 => "11100000",
 5749 => "00011111",
 5750 => "10100110",
 5751 => "10001101",
 5752 => "11011110",
 5753 => "01111111",
 5754 => "00101011",
 5755 => "11011110",
 5756 => "01111010",
 5757 => "00010111",
 5758 => "11100100",
 5759 => "01100010",
 5760 => "10100000",
 5761 => "01010101",
 5762 => "00101111",
 5763 => "10011011",
 5764 => "01011010",
 5765 => "01011111",
 5766 => "00101010",
 5767 => "11001000",
 5768 => "10111100",
 5769 => "10001111",
 5770 => "10111100",
 5771 => "11100110",
 5772 => "10011010",
 5773 => "00001101",
 5774 => "01100101",
 5775 => "01101100",
 5776 => "00100111",
 5777 => "10000110",
 5778 => "10000010",
 5779 => "00011010",
 5780 => "01000100",
 5781 => "00000111",
 5782 => "10110111",
 5783 => "00111000",
 5784 => "11100000",
 5785 => "01011001",
 5786 => "10010011",
 5787 => "01011100",
 5788 => "00100001",
 5789 => "11000111",
 5790 => "10110110",
 5791 => "00011100",
 5792 => "00111100",
 5793 => "11011001",
 5794 => "10110101",
 5795 => "11011001",
 5796 => "01101100",
 5797 => "01001000",
 5798 => "10111101",
 5799 => "10001101",
 5800 => "01011000",
 5801 => "00001100",
 5802 => "10100111",
 5803 => "01011010",
 5804 => "01001100",
 5805 => "11101000",
 5806 => "01001010",
 5807 => "01010010",
 5808 => "01110001",
 5809 => "10111100",
 5810 => "00001011",
 5811 => "11100111",
 5812 => "11110001",
 5813 => "11010110",
 5814 => "01001111",
 5815 => "11010001",
 5816 => "01010101",
 5817 => "01000101",
 5818 => "11100010",
 5819 => "10011010",
 5820 => "00111011",
 5821 => "00100000",
 5822 => "11011110",
 5823 => "10100011",
 5824 => "11010110",
 5825 => "10100000",
 5826 => "10101111",
 5827 => "11110010",
 5828 => "10000011",
 5829 => "01001011",
 5830 => "11011100",
 5831 => "01001100",
 5832 => "00001101",
 5833 => "01111011",
 5834 => "00110001",
 5835 => "10110101",
 5836 => "11011110",
 5837 => "01110110",
 5838 => "00101100",
 5839 => "01001011",
 5840 => "00000101",
 5841 => "01111111",
 5842 => "01100000",
 5843 => "00000010",
 5844 => "01011001",
 5845 => "00101010",
 5846 => "10111011",
 5847 => "11101111",
 5848 => "01101001",
 5849 => "01111011",
 5850 => "01100110",
 5851 => "01101000",
 5852 => "01111011",
 5853 => "10111000",
 5854 => "01110001",
 5855 => "00111001",
 5856 => "10110001",
 5857 => "00010000",
 5858 => "11101000",
 5859 => "00111001",
 5860 => "01111011",
 5861 => "11101011",
 5862 => "11100001",
 5863 => "11011110",
 5864 => "01000100",
 5865 => "10111001",
 5866 => "10111110",
 5867 => "01100010",
 5868 => "01100000",
 5869 => "11111100",
 5870 => "01010011",
 5871 => "01110111",
 5872 => "00001101",
 5873 => "00000111",
 5874 => "11000000",
 5875 => "11101011",
 5876 => "00110001",
 5877 => "10100010",
 5878 => "10101011",
 5879 => "01101011",
 5880 => "01000110",
 5881 => "11001101",
 5882 => "00111100",
 5883 => "00110110",
 5884 => "00010010",
 5885 => "10000010",
 5886 => "01111110",
 5887 => "01111001",
 5888 => "10000101",
 5889 => "00110001",
 5890 => "00011100",
 5891 => "01100001",
 5892 => "01101100",
 5893 => "11101011",
 5894 => "00100001",
 5895 => "00010001",
 5896 => "11101110",
 5897 => "10110000",
 5898 => "00010110",
 5899 => "10111010",
 5900 => "10111100",
 5901 => "00110001",
 5902 => "00000010",
 5903 => "00000011",
 5904 => "11110010",
 5905 => "10010101",
 5906 => "10101110",
 5907 => "10101011",
 5908 => "00000110",
 5909 => "01011101",
 5910 => "10010100",
 5911 => "10001000",
 5912 => "01100011",
 5913 => "10010111",
 5914 => "01101111",
 5915 => "01010000",
 5916 => "00100010",
 5917 => "01000000",
 5918 => "01001000",
 5919 => "00001111",
 5920 => "01100100",
 5921 => "01110000",
 5922 => "01000010",
 5923 => "11010111",
 5924 => "00111001",
 5925 => "11010111",
 5926 => "00011110",
 5927 => "10100110",
 5928 => "10011000",
 5929 => "11011111",
 5930 => "10110000",
 5931 => "10101011",
 5932 => "11000111",
 5933 => "11111111",
 5934 => "10010000",
 5935 => "00011001",
 5936 => "01011011",
 5937 => "10111100",
 5938 => "11101001",
 5939 => "00011010",
 5940 => "01010111",
 5941 => "11101100",
 5942 => "01011101",
 5943 => "11011011",
 5944 => "01101110",
 5945 => "10000100",
 5946 => "00000000",
 5947 => "00110101",
 5948 => "11001010",
 5949 => "00110010",
 5950 => "10111111",
 5951 => "10100101",
 5952 => "11101111",
 5953 => "10011110",
 5954 => "01100011",
 5955 => "11101100",
 5956 => "11101110",
 5957 => "10110010",
 5958 => "11111101",
 5959 => "10001111",
 5960 => "01101011",
 5961 => "00100001",
 5962 => "00001001",
 5963 => "10110110",
 5964 => "11000010",
 5965 => "00010010",
 5966 => "10001111",
 5967 => "01011101",
 5968 => "01011100",
 5969 => "10010110",
 5970 => "10101010",
 5971 => "10000011",
 5972 => "01010001",
 5973 => "10110011",
 5974 => "01001110",
 5975 => "01000101",
 5976 => "01101110",
 5977 => "01111111",
 5978 => "10101000",
 5979 => "00010110",
 5980 => "11110110",
 5981 => "10110110",
 5982 => "01100010",
 5983 => "10100101",
 5984 => "11001000",
 5985 => "10011110",
 5986 => "01011100",
 5987 => "11001010",
 5988 => "01101001",
 5989 => "10100110",
 5990 => "01100110",
 5991 => "00101010",
 5992 => "00100100",
 5993 => "11111010",
 5994 => "01010110",
 5995 => "11011110",
 5996 => "10010010",
 5997 => "10001011",
 5998 => "01011001",
 5999 => "10101111",
 6000 => "11001000",
 6001 => "01110100",
 6002 => "10000001",
 6003 => "10000001",
 6004 => "11011110",
 6005 => "10001011",
 6006 => "00101100",
 6007 => "00001101",
 6008 => "00000001",
 6009 => "11101100",
 6010 => "11001111",
 6011 => "00111011",
 6012 => "01111100",
 6013 => "10110001",
 6014 => "00110100",
 6015 => "00111001",
 6016 => "01111000",
 6017 => "10100110",
 6018 => "11101110",
 6019 => "10001010",
 6020 => "01001100",
 6021 => "11111101",
 6022 => "11011101",
 6023 => "10000110",
 6024 => "11001011",
 6025 => "11111110",
 6026 => "11101111",
 6027 => "11000010",
 6028 => "11011001",
 6029 => "01111001",
 6030 => "01011110",
 6031 => "10000000",
 6032 => "00110101",
 6033 => "11010011",
 6034 => "01110111",
 6035 => "10000110",
 6036 => "01101110",
 6037 => "01111010",
 6038 => "11011010",
 6039 => "00001000",
 6040 => "01101010",
 6041 => "01010011",
 6042 => "10001000",
 6043 => "01111010",
 6044 => "11011110",
 6045 => "00110101",
 6046 => "01001010",
 6047 => "11011011",
 6048 => "10011010",
 6049 => "00110010",
 6050 => "10011000",
 6051 => "01101111",
 6052 => "00010100",
 6053 => "00011110",
 6054 => "01010110",
 6055 => "00011000",
 6056 => "01100111",
 6057 => "11000100",
 6058 => "10000010",
 6059 => "11100010",
 6060 => "11011100",
 6061 => "01000110",
 6062 => "10011001",
 6063 => "01011101",
 6064 => "01010011",
 6065 => "10100110",
 6066 => "00100000",
 6067 => "11101000",
 6068 => "10110100",
 6069 => "11110001",
 6070 => "01111100",
 6071 => "11000011",
 6072 => "10010000",
 6073 => "00011101",
 6074 => "10010111",
 6075 => "00000000",
 6076 => "01110111",
 6077 => "10000110",
 6078 => "00001001",
 6079 => "01000100",
 6080 => "11001001",
 6081 => "01010000",
 6082 => "10100001",
 6083 => "11111110",
 6084 => "00100111",
 6085 => "01000010",
 6086 => "10010100",
 6087 => "11111100",
 6088 => "00100010",
 6089 => "10001011",
 6090 => "00110011",
 6091 => "01100100",
 6092 => "11111111",
 6093 => "01000000",
 6094 => "11100011",
 6095 => "11101101",
 6096 => "11111111",
 6097 => "10010110",
 6098 => "00100000",
 6099 => "00100100",
 6100 => "10010011",
 6101 => "00100010",
 6102 => "11010101",
 6103 => "01100000",
 6104 => "01000010",
 6105 => "10010011",
 6106 => "10110100",
 6107 => "01110110",
 6108 => "00110101",
 6109 => "01101010",
 6110 => "00101100",
 6111 => "00000001",
 6112 => "11110000",
 6113 => "00010100",
 6114 => "11011011",
 6115 => "01100000",
 6116 => "00111110",
 6117 => "01010101",
 6118 => "10010011",
 6119 => "10011101",
 6120 => "10110101",
 6121 => "11111010",
 6122 => "00011000",
 6123 => "10100010",
 6124 => "01001011",
 6125 => "00011010",
 6126 => "10111010",
 6127 => "01010011",
 6128 => "00000100",
 6129 => "10110000",
 6130 => "00100111",
 6131 => "00110110",
 6132 => "00110111",
 6133 => "10100100",
 6134 => "10110100",
 6135 => "00001010",
 6136 => "01100101",
 6137 => "11100000",
 6138 => "01100101",
 6139 => "01000111",
 6140 => "01100101",
 6141 => "10001110",
 6142 => "10110011",
 6143 => "10010100",
 6144 => "10110010",
 6145 => "01111111",
 6146 => "11101111",
 6147 => "11001101",
 6148 => "10010000",
 6149 => "11000100",
 6150 => "00110111",
 6151 => "01110111",
 6152 => "01010010",
 6153 => "00111000",
 6154 => "01011010",
 6155 => "10010000",
 6156 => "11101001",
 6157 => "11101001",
 6158 => "11111100",
 6159 => "11101000",
 6160 => "01001110",
 6161 => "01110000",
 6162 => "10110100",
 6163 => "01000111",
 6164 => "01101101",
 6165 => "11110011",
 6166 => "10001011",
 6167 => "11010100",
 6168 => "10110001",
 6169 => "11110101",
 6170 => "10100111",
 6171 => "11000011",
 6172 => "10001001",
 6173 => "10100111",
 6174 => "10000101",
 6175 => "11100010",
 6176 => "01001000",
 6177 => "10100111",
 6178 => "10110011",
 6179 => "01011100",
 6180 => "11010110",
 6181 => "01110011",
 6182 => "11011010",
 6183 => "10000011",
 6184 => "00000011",
 6185 => "00101011",
 6186 => "10011101",
 6187 => "00110010",
 6188 => "01101001",
 6189 => "11011111",
 6190 => "11011011",
 6191 => "01000001",
 6192 => "00100001",
 6193 => "01100010",
 6194 => "11100101",
 6195 => "01000000",
 6196 => "00111011",
 6197 => "00101110",
 6198 => "00001010",
 6199 => "00100110",
 6200 => "01110000",
 6201 => "00001011",
 6202 => "10101000",
 6203 => "00001100",
 6204 => "01000111",
 6205 => "00000100",
 6206 => "10011010",
 6207 => "11111001",
 6208 => "01010111",
 6209 => "01011010",
 6210 => "11111011",
 6211 => "00010011",
 6212 => "01100100",
 6213 => "11111111",
 6214 => "11111101",
 6215 => "01110011",
 6216 => "10001000",
 6217 => "00111010",
 6218 => "01010101",
 6219 => "00001001",
 6220 => "01011110",
 6221 => "01100100",
 6222 => "01000110",
 6223 => "11000100",
 6224 => "01001000",
 6225 => "01101111",
 6226 => "01110001",
 6227 => "00011100",
 6228 => "11011101",
 6229 => "11110000",
 6230 => "00111101",
 6231 => "01110101",
 6232 => "00010011",
 6233 => "10110100",
 6234 => "10111010",
 6235 => "11001000",
 6236 => "11011111",
 6237 => "01010011",
 6238 => "01111001",
 6239 => "10101111",
 6240 => "10011101",
 6241 => "01111000",
 6242 => "10000111",
 6243 => "11011010",
 6244 => "10010100",
 6245 => "01110011",
 6246 => "11001110",
 6247 => "10011111",
 6248 => "00011111",
 6249 => "11010111",
 6250 => "01101111",
 6251 => "11111110",
 6252 => "10110110",
 6253 => "10010101",
 6254 => "01011100",
 6255 => "01011001",
 6256 => "11100000",
 6257 => "11100001",
 6258 => "11110111",
 6259 => "01011011",
 6260 => "10010111",
 6261 => "00111110",
 6262 => "00101111",
 6263 => "01101110",
 6264 => "00100011",
 6265 => "01010101",
 6266 => "01100010",
 6267 => "11011000",
 6268 => "11010011",
 6269 => "11101111",
 6270 => "01111100",
 6271 => "00110110",
 6272 => "11101100",
 6273 => "11100101",
 6274 => "10101110",
 6275 => "01001011",
 6276 => "00001000",
 6277 => "11000101",
 6278 => "00011011",
 6279 => "01011101",
 6280 => "01110100",
 6281 => "00001101",
 6282 => "00101010",
 6283 => "00000111",
 6284 => "10100111",
 6285 => "00001000",
 6286 => "11100101",
 6287 => "11010101",
 6288 => "01101111",
 6289 => "10111010",
 6290 => "10110101",
 6291 => "01110000",
 6292 => "00110111",
 6293 => "00110101",
 6294 => "10011100",
 6295 => "01111100",
 6296 => "11101011",
 6297 => "01010101",
 6298 => "00100100",
 6299 => "10011010",
 6300 => "11110010",
 6301 => "11110100",
 6302 => "00011010",
 6303 => "10001111",
 6304 => "00001110",
 6305 => "00010010",
 6306 => "10001010",
 6307 => "01111000",
 6308 => "01011011",
 6309 => "11011011",
 6310 => "01110110",
 6311 => "10111110",
 6312 => "01000101",
 6313 => "01101010",
 6314 => "10000010",
 6315 => "11101101",
 6316 => "10111110",
 6317 => "11000010",
 6318 => "01000011",
 6319 => "01000100",
 6320 => "01000110",
 6321 => "00000110",
 6322 => "11010010",
 6323 => "11101111",
 6324 => "00000111",
 6325 => "10000100",
 6326 => "01111111",
 6327 => "10000100",
 6328 => "00110000",
 6329 => "01010101",
 6330 => "01101101",
 6331 => "00011000",
 6332 => "10101010",
 6333 => "01101000",
 6334 => "00000011",
 6335 => "00011100",
 6336 => "01100101",
 6337 => "00010101",
 6338 => "10010001",
 6339 => "10111100",
 6340 => "10001101",
 6341 => "10010010",
 6342 => "10111100",
 6343 => "01001100",
 6344 => "11100101",
 6345 => "00000000",
 6346 => "00001001",
 6347 => "10110110",
 6348 => "01111100",
 6349 => "00110100",
 6350 => "10101000",
 6351 => "10111010",
 6352 => "00010100",
 6353 => "00010011",
 6354 => "01111001",
 6355 => "11010110",
 6356 => "11000011",
 6357 => "11010001",
 6358 => "11100100",
 6359 => "11100101",
 6360 => "11111111",
 6361 => "11111110",
 6362 => "10011001",
 6363 => "10011010",
 6364 => "01011110",
 6365 => "11011100",
 6366 => "01111101",
 6367 => "00010101",
 6368 => "11110000",
 6369 => "01101111",
 6370 => "11010001",
 6371 => "00101100",
 6372 => "10111011",
 6373 => "01010011",
 6374 => "01000110",
 6375 => "00110001",
 6376 => "00101100",
 6377 => "00101111",
 6378 => "01111010",
 6379 => "00011110",
 6380 => "00100001",
 6381 => "10001000",
 6382 => "10011111",
 6383 => "10001001",
 6384 => "10100001",
 6385 => "00000000",
 6386 => "11010100",
 6387 => "00101111",
 6388 => "11101011",
 6389 => "10011101",
 6390 => "11101110",
 6391 => "00101100",
 6392 => "01111000",
 6393 => "01011101",
 6394 => "11010100",
 6395 => "10100010",
 6396 => "01110001",
 6397 => "10001000",
 6398 => "01111101",
 6399 => "10111100",
 6400 => "01110011",
 6401 => "01010000",
 6402 => "11011101",
 6403 => "00000110",
 6404 => "10100101",
 6405 => "00011010",
 6406 => "01100011",
 6407 => "01010110",
 6408 => "00100100",
 6409 => "10110010",
 6410 => "10001101",
 6411 => "10001111",
 6412 => "10011001",
 6413 => "10111110",
 6414 => "11010111",
 6415 => "00110111",
 6416 => "00111001",
 6417 => "00100001",
 6418 => "00000010",
 6419 => "00000111",
 6420 => "00001100",
 6421 => "10110100",
 6422 => "00000110",
 6423 => "11101110",
 6424 => "10011101",
 6425 => "11101100",
 6426 => "10010111",
 6427 => "11101011",
 6428 => "01111100",
 6429 => "11000111",
 6430 => "00110100",
 6431 => "10001111",
 6432 => "11001011",
 6433 => "10001101",
 6434 => "01011001",
 6435 => "11001100",
 6436 => "01111010",
 6437 => "01100111",
 6438 => "01111000",
 6439 => "01110000",
 6440 => "00000100",
 6441 => "11111001",
 6442 => "00011010",
 6443 => "00000111",
 6444 => "01111101",
 6445 => "01100101",
 6446 => "11101101",
 6447 => "11011000",
 6448 => "01100101",
 6449 => "10100111",
 6450 => "10111011",
 6451 => "01010011",
 6452 => "01110011",
 6453 => "00101001",
 6454 => "01000010",
 6455 => "01100101",
 6456 => "00111111",
 6457 => "10000110",
 6458 => "01011001",
 6459 => "01101110",
 6460 => "10111011",
 6461 => "10011010",
 6462 => "10011000",
 6463 => "01010110",
 6464 => "11101010",
 6465 => "01000100",
 6466 => "11001000",
 6467 => "10110110",
 6468 => "01111100",
 6469 => "10000000",
 6470 => "10100101",
 6471 => "10011110",
 6472 => "00010011",
 6473 => "01111011",
 6474 => "00011010",
 6475 => "10100111",
 6476 => "10101001",
 6477 => "11110010",
 6478 => "11111110",
 6479 => "01000010",
 6480 => "01111000",
 6481 => "01000101",
 6482 => "11100101",
 6483 => "11100010",
 6484 => "11001000",
 6485 => "00001011",
 6486 => "11110010",
 6487 => "10111100",
 6488 => "10110000",
 6489 => "00110100",
 6490 => "01000010",
 6491 => "11001100",
 6492 => "01101000",
 6493 => "10010010",
 6494 => "01100011",
 6495 => "11010011",
 6496 => "00101110",
 6497 => "01010101",
 6498 => "11001011",
 6499 => "01010101",
 6500 => "01011101",
 6501 => "00110110",
 6502 => "00001001",
 6503 => "01111110",
 6504 => "10111110",
 6505 => "10110110",
 6506 => "01100110",
 6507 => "11110001",
 6508 => "10011001",
 6509 => "11011011",
 6510 => "00000010",
 6511 => "01101100",
 6512 => "10010000",
 6513 => "11111011",
 6514 => "10101000",
 6515 => "11110010",
 6516 => "01111101",
 6517 => "11100100",
 6518 => "10100110",
 6519 => "00111001",
 6520 => "00101110",
 6521 => "10100000",
 6522 => "10000001",
 6523 => "01001001",
 6524 => "00001100",
 6525 => "00001011",
 6526 => "01001111",
 6527 => "11101101",
 6528 => "11011100",
 6529 => "01010011",
 6530 => "01010000",
 6531 => "00011010",
 6532 => "10111010",
 6533 => "10100010",
 6534 => "01001101",
 6535 => "10100100",
 6536 => "11010111",
 6537 => "00101101",
 6538 => "10011100",
 6539 => "10001011",
 6540 => "10111001",
 6541 => "10101111",
 6542 => "00100101",
 6543 => "00010101",
 6544 => "10100100",
 6545 => "01000100",
 6546 => "00111111",
 6547 => "11001110",
 6548 => "11110000",
 6549 => "00111110",
 6550 => "01010100",
 6551 => "11000101",
 6552 => "10000100",
 6553 => "10100111",
 6554 => "10010111",
 6555 => "00001011",
 6556 => "01101001",
 6557 => "01100110",
 6558 => "01010001",
 6559 => "00010110",
 6560 => "01010100",
 6561 => "01011001",
 6562 => "00100111",
 6563 => "11111010",
 6564 => "01010011",
 6565 => "10001100",
 6566 => "01100011",
 6567 => "00010110",
 6568 => "01101100",
 6569 => "00001101",
 6570 => "00100011",
 6571 => "11110100",
 6572 => "11010010",
 6573 => "11101011",
 6574 => "11011100",
 6575 => "00110111",
 6576 => "11110111",
 6577 => "10010111",
 6578 => "00101000",
 6579 => "10011001",
 6580 => "11101011",
 6581 => "11011010",
 6582 => "11010000",
 6583 => "00111010",
 6584 => "01001100",
 6585 => "11111011",
 6586 => "10111111",
 6587 => "11011000",
 6588 => "10100100",
 6589 => "11000010",
 6590 => "01110000",
 6591 => "10101010",
 6592 => "00100010",
 6593 => "11001000",
 6594 => "10111010",
 6595 => "00011000",
 6596 => "00101000",
 6597 => "11111001",
 6598 => "11110101",
 6599 => "00011111",
 6600 => "10111111",
 6601 => "00010011",
 6602 => "10011011",
 6603 => "00001011",
 6604 => "11000001",
 6605 => "01010111",
 6606 => "10011101",
 6607 => "00011110",
 6608 => "01001011",
 6609 => "01100010",
 6610 => "00100100",
 6611 => "01111111",
 6612 => "11101110",
 6613 => "01101101",
 6614 => "11100000",
 6615 => "10001001",
 6616 => "10110000",
 6617 => "10011101",
 6618 => "00100011",
 6619 => "00110011",
 6620 => "10000101",
 6621 => "00000110",
 6622 => "11001010",
 6623 => "00010011",
 6624 => "11001100",
 6625 => "00001000",
 6626 => "01100011",
 6627 => "10001000",
 6628 => "10001000",
 6629 => "01110100",
 6630 => "01100100",
 6631 => "11000101",
 6632 => "00111011",
 6633 => "01111110",
 6634 => "11111100",
 6635 => "00001110",
 6636 => "00001110",
 6637 => "10101010",
 6638 => "10001101",
 6639 => "00110110",
 6640 => "00100000",
 6641 => "01010001",
 6642 => "10100000",
 6643 => "01110100",
 6644 => "01100110",
 6645 => "10010101",
 6646 => "00011111",
 6647 => "00000101",
 6648 => "11101111",
 6649 => "10100110",
 6650 => "10110101",
 6651 => "11110111",
 6652 => "10010010",
 6653 => "11101100",
 6654 => "01110000",
 6655 => "00000100",
 6656 => "01101001",
 6657 => "10000000",
 6658 => "00100100",
 6659 => "10101111",
 6660 => "10010100",
 6661 => "00111011",
 6662 => "10011111",
 6663 => "11011101",
 6664 => "01101111",
 6665 => "00100000",
 6666 => "11100101",
 6667 => "00110110",
 6668 => "11111110",
 6669 => "01100010",
 6670 => "00100111",
 6671 => "01111011",
 6672 => "10000000",
 6673 => "00010101",
 6674 => "00100110",
 6675 => "00010101",
 6676 => "11001110",
 6677 => "11010111",
 6678 => "00010010",
 6679 => "01111010",
 6680 => "01101110",
 6681 => "10101101",
 6682 => "11110110",
 6683 => "11000100",
 6684 => "00110111",
 6685 => "01110010",
 6686 => "10101001",
 6687 => "00001111",
 6688 => "00101100",
 6689 => "00111011",
 6690 => "10010111",
 6691 => "00110101",
 6692 => "10000011",
 6693 => "00000111",
 6694 => "11000001",
 6695 => "01001001",
 6696 => "10101111",
 6697 => "01101101",
 6698 => "10110111",
 6699 => "10110100",
 6700 => "00111000",
 6701 => "11010101",
 6702 => "10010101",
 6703 => "10000101",
 6704 => "10001001",
 6705 => "10101101",
 6706 => "00001000",
 6707 => "11110100",
 6708 => "00111100",
 6709 => "10010101",
 6710 => "00100001",
 6711 => "11111110",
 6712 => "01110100",
 6713 => "11110001",
 6714 => "10111000",
 6715 => "11001010",
 6716 => "11010000",
 6717 => "11111010",
 6718 => "11110101",
 6719 => "01101111",
 6720 => "01000101",
 6721 => "00100101",
 6722 => "11001010",
 6723 => "01110011",
 6724 => "10001101",
 6725 => "00100100",
 6726 => "00111101",
 6727 => "11011011",
 6728 => "10011010",
 6729 => "00011101",
 6730 => "11010101",
 6731 => "00010111",
 6732 => "11101111",
 6733 => "10010011",
 6734 => "01010011",
 6735 => "10000010",
 6736 => "00010000",
 6737 => "00101101",
 6738 => "01110011",
 6739 => "10111101",
 6740 => "00111110",
 6741 => "01010111",
 6742 => "11110000",
 6743 => "11110100",
 6744 => "10101111",
 6745 => "00110001",
 6746 => "10111010",
 6747 => "01110000",
 6748 => "00011101",
 6749 => "00011000",
 6750 => "01001111",
 6751 => "10000111",
 6752 => "11101001",
 6753 => "00100100",
 6754 => "00101101",
 6755 => "10011100",
 6756 => "10000001",
 6757 => "01010000",
 6758 => "10110001",
 6759 => "00100001",
 6760 => "00100111",
 6761 => "01111100",
 6762 => "01110110",
 6763 => "10010011",
 6764 => "00001010",
 6765 => "11100100",
 6766 => "10000100",
 6767 => "00100000",
 6768 => "00111000",
 6769 => "00100100",
 6770 => "01110110",
 6771 => "00101001",
 6772 => "11100000",
 6773 => "10110100",
 6774 => "10010001",
 6775 => "01101111",
 6776 => "01110000",
 6777 => "01101000",
 6778 => "10111111",
 6779 => "10010000",
 6780 => "11101000",
 6781 => "01101001",
 6782 => "01100110",
 6783 => "00001100",
 6784 => "00110000",
 6785 => "11010100",
 6786 => "00111110",
 6787 => "11000000",
 6788 => "10000010",
 6789 => "11111000",
 6790 => "00111100",
 6791 => "01000111",
 6792 => "01000110",
 6793 => "11001110",
 6794 => "10111110",
 6795 => "01011110",
 6796 => "10100110",
 6797 => "01110010",
 6798 => "01010111",
 6799 => "11111011",
 6800 => "11011011",
 6801 => "01100100",
 6802 => "00110111",
 6803 => "11011101",
 6804 => "11111110",
 6805 => "01010000",
 6806 => "10000000",
 6807 => "10111011",
 6808 => "00110011",
 6809 => "01011011",
 6810 => "10000000",
 6811 => "01011011",
 6812 => "11101011",
 6813 => "01000001",
 6814 => "01001000",
 6815 => "00011010",
 6816 => "00101101",
 6817 => "10110001",
 6818 => "11000010",
 6819 => "11011011",
 6820 => "00001110",
 6821 => "01100100",
 6822 => "01010000",
 6823 => "01110000",
 6824 => "01111100",
 6825 => "00001011",
 6826 => "01000100",
 6827 => "10100100",
 6828 => "00100000",
 6829 => "00001000",
 6830 => "01001011",
 6831 => "01001100",
 6832 => "10011110",
 6833 => "10111100",
 6834 => "10000001",
 6835 => "11101111",
 6836 => "00001000",
 6837 => "01100011",
 6838 => "00011001",
 6839 => "00011000",
 6840 => "10000111",
 6841 => "01100011",
 6842 => "10100000",
 6843 => "01000000",
 6844 => "01100110",
 6845 => "11000001",
 6846 => "10101011",
 6847 => "01100001",
 6848 => "00100011",
 6849 => "10100010",
 6850 => "01001011",
 6851 => "11010010",
 6852 => "01011111",
 6853 => "11101001",
 6854 => "11100111",
 6855 => "01111001",
 6856 => "01110101",
 6857 => "01001010",
 6858 => "10111011",
 6859 => "11001110",
 6860 => "01010010",
 6861 => "01111100",
 6862 => "00000111",
 6863 => "00110101",
 6864 => "10100100",
 6865 => "11000111",
 6866 => "00101011",
 6867 => "01101100",
 6868 => "10001101",
 6869 => "11110010",
 6870 => "11100000",
 6871 => "00001001",
 6872 => "01100110",
 6873 => "11111110",
 6874 => "11010010",
 6875 => "10000001",
 6876 => "11110000",
 6877 => "10111111",
 6878 => "01010000",
 6879 => "10111001",
 6880 => "01101100",
 6881 => "10011100",
 6882 => "11100101",
 6883 => "00101100",
 6884 => "10001010",
 6885 => "10110110",
 6886 => "11111101",
 6887 => "01011001",
 6888 => "11101100",
 6889 => "01000000",
 6890 => "00010101",
 6891 => "11011010",
 6892 => "00110010",
 6893 => "10110010",
 6894 => "11011110",
 6895 => "01110100",
 6896 => "11111011",
 6897 => "11110001",
 6898 => "01001111",
 6899 => "00001010",
 6900 => "11100110",
 6901 => "11110001",
 6902 => "10101010",
 6903 => "00100101",
 6904 => "00011010",
 6905 => "00000001",
 6906 => "11001111",
 6907 => "11100100",
 6908 => "00110010",
 6909 => "01110100",
 6910 => "11110011",
 6911 => "00101000",
 6912 => "11000010",
 6913 => "01110000",
 6914 => "00100100",
 6915 => "01011001",
 6916 => "00100010",
 6917 => "00100010",
 6918 => "11011100",
 6919 => "01010111",
 6920 => "00011111",
 6921 => "11000010",
 6922 => "01011110",
 6923 => "10000100",
 6924 => "10111101",
 6925 => "01111001",
 6926 => "11111011",
 6927 => "00010111",
 6928 => "11000110",
 6929 => "11010100",
 6930 => "10101100",
 6931 => "00110000",
 6932 => "01100111",
 6933 => "11110000",
 6934 => "10100001",
 6935 => "01011100",
 6936 => "11100010",
 6937 => "11101000",
 6938 => "11100011",
 6939 => "10111001",
 6940 => "00100011",
 6941 => "01000110",
 6942 => "11110111",
 6943 => "11011011",
 6944 => "01111011",
 6945 => "11100001",
 6946 => "01111111",
 6947 => "00101010",
 6948 => "01110111",
 6949 => "11100000",
 6950 => "01000101",
 6951 => "01001011",
 6952 => "11111010",
 6953 => "00101101",
 6954 => "00000001",
 6955 => "00001101",
 6956 => "10111010",
 6957 => "10011010",
 6958 => "11111100",
 6959 => "00011111",
 6960 => "10011001",
 6961 => "11111111",
 6962 => "10101010",
 6963 => "11010100",
 6964 => "01111011",
 6965 => "01101000",
 6966 => "01011111",
 6967 => "01010011",
 6968 => "11100100",
 6969 => "01100110",
 6970 => "01100011",
 6971 => "11101011",
 6972 => "11111011",
 6973 => "10111001",
 6974 => "00010110",
 6975 => "11111100",
 6976 => "10000011",
 6977 => "01111001",
 6978 => "10110101",
 6979 => "00100111",
 6980 => "10111111",
 6981 => "01001111",
 6982 => "10001010",
 6983 => "01110000",
 6984 => "00111111",
 6985 => "10100010",
 6986 => "01000011",
 6987 => "11000101",
 6988 => "10010101",
 6989 => "01010010",
 6990 => "01010011",
 6991 => "11000011",
 6992 => "11000001",
 6993 => "10110010",
 6994 => "10100011",
 6995 => "01101000",
 6996 => "01110011",
 6997 => "00111110",
 6998 => "11001100",
 6999 => "00111001",
 7000 => "10000001",
 7001 => "10001010",
 7002 => "00110110",
 7003 => "01001101",
 7004 => "10111010",
 7005 => "10001000",
 7006 => "11000111",
 7007 => "01000111",
 7008 => "01001011",
 7009 => "00000101",
 7010 => "01011100",
 7011 => "11101110",
 7012 => "00110110",
 7013 => "00001011",
 7014 => "11010010",
 7015 => "11001000",
 7016 => "01001000",
 7017 => "00110101",
 7018 => "10010010",
 7019 => "00000000",
 7020 => "10000100",
 7021 => "11110000",
 7022 => "01110001",
 7023 => "01100010",
 7024 => "11011110",
 7025 => "11101011",
 7026 => "10001100",
 7027 => "01001101",
 7028 => "10101110",
 7029 => "10011101",
 7030 => "01001110",
 7031 => "10001001",
 7032 => "11011101",
 7033 => "11000101",
 7034 => "00001110",
 7035 => "10001010",
 7036 => "11110010",
 7037 => "10001101",
 7038 => "10101001",
 7039 => "11001011",
 7040 => "01001101",
 7041 => "10111101",
 7042 => "01010100",
 7043 => "00110010",
 7044 => "10100000",
 7045 => "00111011",
 7046 => "11001111",
 7047 => "10001101",
 7048 => "00110011",
 7049 => "11110101",
 7050 => "11000110",
 7051 => "00010101",
 7052 => "01110100",
 7053 => "00100011",
 7054 => "01010111",
 7055 => "01110001",
 7056 => "00011101",
 7057 => "10100100",
 7058 => "01101000",
 7059 => "01010010",
 7060 => "01010111",
 7061 => "11100011",
 7062 => "01010110",
 7063 => "11100111",
 7064 => "11001101",
 7065 => "11011110",
 7066 => "01100011",
 7067 => "00010001",
 7068 => "10011001",
 7069 => "01110101",
 7070 => "11110100",
 7071 => "11001100",
 7072 => "00011010",
 7073 => "11010000",
 7074 => "10010101",
 7075 => "00011011",
 7076 => "00001001",
 7077 => "10010100",
 7078 => "00110011",
 7079 => "01011011",
 7080 => "01011010",
 7081 => "00101100",
 7082 => "01010001",
 7083 => "11110110",
 7084 => "11000010",
 7085 => "10001101",
 7086 => "01011011",
 7087 => "00011011",
 7088 => "10111100",
 7089 => "10100101",
 7090 => "11110100",
 7091 => "11011011",
 7092 => "11110100",
 7093 => "11101111",
 7094 => "00111111",
 7095 => "10100000",
 7096 => "11100011",
 7097 => "00001110",
 7098 => "11011110",
 7099 => "01011010",
 7100 => "01101111",
 7101 => "10010001",
 7102 => "01001110",
 7103 => "11100110",
 7104 => "10000100",
 7105 => "00110001",
 7106 => "11000111",
 7107 => "11001011",
 7108 => "11111110",
 7109 => "00100010",
 7110 => "11111110",
 7111 => "10000100",
 7112 => "10111000",
 7113 => "00000010",
 7114 => "11000110",
 7115 => "11111010",
 7116 => "00000110",
 7117 => "01010101",
 7118 => "00100110",
 7119 => "01001000",
 7120 => "11010110",
 7121 => "11001101",
 7122 => "10010110",
 7123 => "01010100",
 7124 => "01101101",
 7125 => "10001111",
 7126 => "11000000",
 7127 => "00100010",
 7128 => "01101101",
 7129 => "10000011",
 7130 => "10001111",
 7131 => "10101101",
 7132 => "00110111",
 7133 => "01000010",
 7134 => "01110111",
 7135 => "00100101",
 7136 => "10011011",
 7137 => "10100001",
 7138 => "01000111",
 7139 => "01101001",
 7140 => "00010001",
 7141 => "11110100",
 7142 => "10110000",
 7143 => "01101111",
 7144 => "10000000",
 7145 => "00000110",
 7146 => "01101000",
 7147 => "00011110",
 7148 => "10000100",
 7149 => "10111110",
 7150 => "10111100",
 7151 => "00111001",
 7152 => "11110110",
 7153 => "11110010",
 7154 => "11101000",
 7155 => "11100010",
 7156 => "11001000",
 7157 => "00101000",
 7158 => "00101011",
 7159 => "00010011",
 7160 => "10010010",
 7161 => "01011001",
 7162 => "00110010",
 7163 => "10000000",
 7164 => "00011011",
 7165 => "11100111",
 7166 => "01111010",
 7167 => "11111000",
 7168 => "11010111",
 7169 => "11100000",
 7170 => "01111010",
 7171 => "10010000",
 7172 => "01010110",
 7173 => "10110000",
 7174 => "11000101",
 7175 => "01000100",
 7176 => "01000010",
 7177 => "11001010",
 7178 => "00001111",
 7179 => "10001100",
 7180 => "11000011",
 7181 => "10000111",
 7182 => "01010101",
 7183 => "10010101",
 7184 => "00000110",
 7185 => "11001110",
 7186 => "00011111",
 7187 => "11010011",
 7188 => "00001110",
 7189 => "10001000",
 7190 => "10101111",
 7191 => "00011010",
 7192 => "11111000",
 7193 => "10101101",
 7194 => "10100100",
 7195 => "11010001",
 7196 => "00011011",
 7197 => "01001111",
 7198 => "11111001",
 7199 => "00111001",
 7200 => "01001101",
 7201 => "11011111",
 7202 => "11011101",
 7203 => "00100010",
 7204 => "11000110",
 7205 => "01100100",
 7206 => "11101010",
 7207 => "11100110",
 7208 => "10110110",
 7209 => "00001111",
 7210 => "10100101",
 7211 => "11101110",
 7212 => "10100010",
 7213 => "10111110",
 7214 => "10100100",
 7215 => "00111010",
 7216 => "01011110",
 7217 => "00010011",
 7218 => "11000110",
 7219 => "11101111",
 7220 => "11110111",
 7221 => "00101101",
 7222 => "10110110",
 7223 => "10001100",
 7224 => "10110011",
 7225 => "10101100",
 7226 => "10010100",
 7227 => "01111001",
 7228 => "10011010",
 7229 => "00111110",
 7230 => "11010000",
 7231 => "11101111",
 7232 => "01011011",
 7233 => "00011111",
 7234 => "11010000",
 7235 => "11011110",
 7236 => "01100110",
 7237 => "01110001",
 7238 => "10111110",
 7239 => "00000011",
 7240 => "10101100",
 7241 => "10110010",
 7242 => "11011100",
 7243 => "11011101",
 7244 => "01000100",
 7245 => "00011100",
 7246 => "01101001",
 7247 => "10000111",
 7248 => "11000001",
 7249 => "11101111",
 7250 => "10101001",
 7251 => "00001111",
 7252 => "11010001",
 7253 => "00001010",
 7254 => "11111000",
 7255 => "11101101",
 7256 => "00010000",
 7257 => "01100101",
 7258 => "10110101",
 7259 => "01110001",
 7260 => "11110101",
 7261 => "00110111",
 7262 => "01101001",
 7263 => "10010111",
 7264 => "00000101",
 7265 => "00011011",
 7266 => "00010100",
 7267 => "11111000",
 7268 => "00111111",
 7269 => "01010000",
 7270 => "00011111",
 7271 => "01010000",
 7272 => "01000011",
 7273 => "01001011",
 7274 => "00101001",
 7275 => "10100110",
 7276 => "00001101",
 7277 => "10111001",
 7278 => "00111001",
 7279 => "01010100",
 7280 => "01100010",
 7281 => "00111001",
 7282 => "00110111",
 7283 => "10000110",
 7284 => "11110100",
 7285 => "10000101",
 7286 => "10010110",
 7287 => "11101110",
 7288 => "10010000",
 7289 => "10001101",
 7290 => "00100110",
 7291 => "00100010",
 7292 => "01111000",
 7293 => "11111011",
 7294 => "10101011",
 7295 => "10111111",
 7296 => "00101110",
 7297 => "01010101",
 7298 => "00001001",
 7299 => "11000000",
 7300 => "11110101",
 7301 => "10100111",
 7302 => "10001011",
 7303 => "00010000",
 7304 => "11111110",
 7305 => "11100100",
 7306 => "01010100",
 7307 => "00001010",
 7308 => "10000100",
 7309 => "01011010",
 7310 => "11111101",
 7311 => "00010111",
 7312 => "01011100",
 7313 => "00001000",
 7314 => "01011100",
 7315 => "00011010",
 7316 => "10010000",
 7317 => "10010110",
 7318 => "11100010",
 7319 => "00100111",
 7320 => "00010000",
 7321 => "11110110",
 7322 => "10101101",
 7323 => "11100000",
 7324 => "00001011",
 7325 => "11101100",
 7326 => "11011001",
 7327 => "11111010",
 7328 => "11111100",
 7329 => "01111111",
 7330 => "01000100",
 7331 => "00100110",
 7332 => "01000001",
 7333 => "11111101",
 7334 => "00101011",
 7335 => "01011000",
 7336 => "01110011",
 7337 => "01101001",
 7338 => "01100010",
 7339 => "10011000",
 7340 => "00110011",
 7341 => "11101101",
 7342 => "01000001",
 7343 => "00110000",
 7344 => "10001110",
 7345 => "01100101",
 7346 => "11001111",
 7347 => "11011000",
 7348 => "01000000",
 7349 => "11110001",
 7350 => "11100011",
 7351 => "11111100",
 7352 => "00110111",
 7353 => "10011110",
 7354 => "01100101",
 7355 => "01001100",
 7356 => "11100011",
 7357 => "11111010",
 7358 => "00010000",
 7359 => "10010000",
 7360 => "11100110",
 7361 => "11010101",
 7362 => "11101101",
 7363 => "00000000",
 7364 => "10001100",
 7365 => "00100010",
 7366 => "11010010",
 7367 => "01010011",
 7368 => "01000110",
 7369 => "01101101",
 7370 => "00110010",
 7371 => "00110110",
 7372 => "11011001",
 7373 => "00011111",
 7374 => "01101001",
 7375 => "00001110",
 7376 => "00010000",
 7377 => "10111010",
 7378 => "11000011",
 7379 => "00100111",
 7380 => "11100011",
 7381 => "00100100",
 7382 => "01000011",
 7383 => "10110010",
 7384 => "10010101",
 7385 => "00111111",
 7386 => "00001010",
 7387 => "11010010",
 7388 => "01111111",
 7389 => "00001101",
 7390 => "10010110",
 7391 => "11111011",
 7392 => "00011011",
 7393 => "10101110",
 7394 => "11011101",
 7395 => "00100001",
 7396 => "01011101",
 7397 => "00010111",
 7398 => "11000101",
 7399 => "11100100",
 7400 => "00010011",
 7401 => "01001101",
 7402 => "10100010",
 7403 => "11111000",
 7404 => "00100101",
 7405 => "11011100",
 7406 => "01110010",
 7407 => "11001010",
 7408 => "11110001",
 7409 => "10110011",
 7410 => "00010100",
 7411 => "01111101",
 7412 => "10011100",
 7413 => "10010111",
 7414 => "10000001",
 7415 => "11000001",
 7416 => "10011101",
 7417 => "10100110",
 7418 => "10010101",
 7419 => "00000101",
 7420 => "01001010",
 7421 => "11011000",
 7422 => "00111000",
 7423 => "10100001",
 7424 => "00100100",
 7425 => "01111010",
 7426 => "01110011",
 7427 => "10010100",
 7428 => "11100000",
 7429 => "11000110",
 7430 => "01101100",
 7431 => "00111010",
 7432 => "10001001",
 7433 => "10001011",
 7434 => "10000001",
 7435 => "11100001",
 7436 => "11101001",
 7437 => "11101000",
 7438 => "10000010",
 7439 => "11001011",
 7440 => "11010100",
 7441 => "01011110",
 7442 => "11000100",
 7443 => "11101101",
 7444 => "11000100",
 7445 => "01111000",
 7446 => "00000001",
 7447 => "00010001",
 7448 => "10110000",
 7449 => "11101101",
 7450 => "01001011",
 7451 => "01111010",
 7452 => "10110110",
 7453 => "00001011",
 7454 => "00111010",
 7455 => "10110101",
 7456 => "00011010",
 7457 => "10100110",
 7458 => "11010001",
 7459 => "01001111",
 7460 => "11010010",
 7461 => "10110111",
 7462 => "00001001",
 7463 => "01010110",
 7464 => "01001010",
 7465 => "10010001",
 7466 => "10000001",
 7467 => "10110110",
 7468 => "01101010",
 7469 => "11100111",
 7470 => "01110100",
 7471 => "11111111",
 7472 => "00101000",
 7473 => "10100101",
 7474 => "10101000",
 7475 => "01110110",
 7476 => "01111101",
 7477 => "01000101",
 7478 => "10101110",
 7479 => "11010010",
 7480 => "01100111",
 7481 => "00101000",
 7482 => "00000011",
 7483 => "00100110",
 7484 => "01011000",
 7485 => "11110110",
 7486 => "00101010",
 7487 => "11110001",
 7488 => "01001111",
 7489 => "11010100",
 7490 => "01011111",
 7491 => "01000011",
 7492 => "10001011",
 7493 => "11011010",
 7494 => "10001000",
 7495 => "00010000",
 7496 => "01011100",
 7497 => "00111100",
 7498 => "01001101",
 7499 => "10001000",
 7500 => "00000100",
 7501 => "11010100",
 7502 => "01101011",
 7503 => "01001010",
 7504 => "01110100",
 7505 => "01111111",
 7506 => "00010111",
 7507 => "01100100",
 7508 => "01001000",
 7509 => "11111010",
 7510 => "11010011",
 7511 => "11001010",
 7512 => "11010100",
 7513 => "11110111",
 7514 => "10100010",
 7515 => "00001100",
 7516 => "00101110",
 7517 => "01001011",
 7518 => "11011011",
 7519 => "10110111",
 7520 => "00010010",
 7521 => "00111010",
 7522 => "00101101",
 7523 => "01101100",
 7524 => "11000010",
 7525 => "11111010",
 7526 => "00000101",
 7527 => "11010001",
 7528 => "10111110",
 7529 => "10011110",
 7530 => "01010011",
 7531 => "11000010",
 7532 => "11100111",
 7533 => "01111101",
 7534 => "00000001",
 7535 => "00000001",
 7536 => "00000010",
 7537 => "11011100",
 7538 => "01101001",
 7539 => "00111100",
 7540 => "11110010",
 7541 => "01100000",
 7542 => "01111101",
 7543 => "10101000",
 7544 => "11010100",
 7545 => "01110001",
 7546 => "01100100",
 7547 => "00111000",
 7548 => "01000001",
 7549 => "10001100",
 7550 => "00000000",
 7551 => "11111110",
 7552 => "11000111",
 7553 => "10011011",
 7554 => "11010011",
 7555 => "11010001",
 7556 => "11110010",
 7557 => "00111101",
 7558 => "01111001",
 7559 => "01100001",
 7560 => "11010000",
 7561 => "10011111",
 7562 => "01000001",
 7563 => "00000011",
 7564 => "01011110",
 7565 => "00111001",
 7566 => "00101110",
 7567 => "11100100",
 7568 => "10111010",
 7569 => "10001010",
 7570 => "00000100",
 7571 => "11010001",
 7572 => "01001110",
 7573 => "11001000",
 7574 => "00010100",
 7575 => "01100000",
 7576 => "10111001",
 7577 => "10001101",
 7578 => "11100110",
 7579 => "10000100",
 7580 => "10110111",
 7581 => "01101000",
 7582 => "00011011",
 7583 => "01110110",
 7584 => "01101000",
 7585 => "11011100",
 7586 => "11010011",
 7587 => "10011010",
 7588 => "00000000",
 7589 => "10100101",
 7590 => "00010110",
 7591 => "00100010",
 7592 => "01000110",
 7593 => "11001101",
 7594 => "00000000",
 7595 => "10010001",
 7596 => "11011010",
 7597 => "00000011",
 7598 => "10010110",
 7599 => "00111101",
 7600 => "01011101",
 7601 => "00100000",
 7602 => "00100000",
 7603 => "00101001",
 7604 => "00000100",
 7605 => "01010100",
 7606 => "10000101",
 7607 => "00101101",
 7608 => "11101101",
 7609 => "10000011",
 7610 => "01001100",
 7611 => "10111101",
 7612 => "00111100",
 7613 => "00001011",
 7614 => "01000111",
 7615 => "00000001",
 7616 => "01011011",
 7617 => "00100011",
 7618 => "11111011",
 7619 => "10111100",
 7620 => "00100100",
 7621 => "01010101",
 7622 => "01001101",
 7623 => "01111110",
 7624 => "11001010",
 7625 => "00001111",
 7626 => "11100100",
 7627 => "11111010",
 7628 => "11000001",
 7629 => "10111010",
 7630 => "00000101",
 7631 => "11111001",
 7632 => "11111111",
 7633 => "01111110",
 7634 => "00011101",
 7635 => "00100000",
 7636 => "01010000",
 7637 => "01000001",
 7638 => "00011000",
 7639 => "01010110",
 7640 => "01011101",
 7641 => "00110110",
 7642 => "01001000",
 7643 => "10011100",
 7644 => "10001010",
 7645 => "11100000",
 7646 => "01011110",
 7647 => "01001100",
 7648 => "10000111",
 7649 => "01011000",
 7650 => "00000111",
 7651 => "10011001",
 7652 => "10101110",
 7653 => "01001101",
 7654 => "10111001",
 7655 => "11001000",
 7656 => "10101101",
 7657 => "10111000",
 7658 => "00010000",
 7659 => "00100111",
 7660 => "01000010",
 7661 => "10011001",
 7662 => "11011101",
 7663 => "00110010",
 7664 => "10001011",
 7665 => "00000110",
 7666 => "11001100",
 7667 => "01111111",
 7668 => "11001000",
 7669 => "01101110",
 7670 => "11010011",
 7671 => "00010000",
 7672 => "01011000",
 7673 => "10001001",
 7674 => "00010010",
 7675 => "10011001",
 7676 => "10000011",
 7677 => "10001010",
 7678 => "11100100",
 7679 => "01001111",
 7680 => "11111011",
 7681 => "11100111",
 7682 => "10011111",
 7683 => "01110010",
 7684 => "11001111",
 7685 => "01000011",
 7686 => "01101100",
 7687 => "00011111",
 7688 => "01000110",
 7689 => "00111010",
 7690 => "00000101",
 7691 => "00000111",
 7692 => "00101100",
 7693 => "01110110",
 7694 => "10001011",
 7695 => "00010001",
 7696 => "01111111",
 7697 => "01111010",
 7698 => "00011000",
 7699 => "01010011",
 7700 => "11010011",
 7701 => "10011001",
 7702 => "00011100",
 7703 => "11111100",
 7704 => "00101100",
 7705 => "00001111",
 7706 => "11110100",
 7707 => "10111001",
 7708 => "01010011",
 7709 => "00111010",
 7710 => "11010001",
 7711 => "10010011",
 7712 => "10101101",
 7713 => "11001011",
 7714 => "01111111",
 7715 => "00000111",
 7716 => "00100000",
 7717 => "01010111",
 7718 => "01100010",
 7719 => "01000100",
 7720 => "00111101",
 7721 => "10111101",
 7722 => "11010111",
 7723 => "01111110",
 7724 => "00100110",
 7725 => "01001100",
 7726 => "10111000",
 7727 => "01110011",
 7728 => "10101101",
 7729 => "11011100",
 7730 => "00110011",
 7731 => "00101001",
 7732 => "11111001",
 7733 => "11101010",
 7734 => "11100100",
 7735 => "11000111",
 7736 => "01000010",
 7737 => "01100000",
 7738 => "11101000",
 7739 => "11101010",
 7740 => "10111000",
 7741 => "11100110",
 7742 => "11101000",
 7743 => "10101001",
 7744 => "10100111",
 7745 => "00011100",
 7746 => "10000001",
 7747 => "10100100",
 7748 => "10110001",
 7749 => "00001100",
 7750 => "11101110",
 7751 => "01100101",
 7752 => "01111001",
 7753 => "10111100",
 7754 => "10011000",
 7755 => "10110111",
 7756 => "01111101",
 7757 => "01010101",
 7758 => "01111001",
 7759 => "10101010",
 7760 => "00000100",
 7761 => "11100100",
 7762 => "01010001",
 7763 => "01000100",
 7764 => "01111011",
 7765 => "00010011",
 7766 => "11110000",
 7767 => "01011001",
 7768 => "11101110",
 7769 => "10011000",
 7770 => "10011110",
 7771 => "11111001",
 7772 => "00100010",
 7773 => "10000010",
 7774 => "10110001",
 7775 => "11010001",
 7776 => "11000010",
 7777 => "00011101",
 7778 => "00110010",
 7779 => "11001100",
 7780 => "01100011",
 7781 => "01111110",
 7782 => "10000000",
 7783 => "00110001",
 7784 => "00010011",
 7785 => "01110000",
 7786 => "11001101",
 7787 => "10101110",
 7788 => "01011101",
 7789 => "01100011",
 7790 => "00011111",
 7791 => "00001010",
 7792 => "11100110",
 7793 => "01001001",
 7794 => "11010101",
 7795 => "11110011",
 7796 => "10110000",
 7797 => "00011011",
 7798 => "00110101",
 7799 => "11110100",
 7800 => "00110011",
 7801 => "01111011",
 7802 => "10010100",
 7803 => "00000011",
 7804 => "01110010",
 7805 => "01101100",
 7806 => "00011101",
 7807 => "01111011",
 7808 => "11111001",
 7809 => "00011110",
 7810 => "11011101",
 7811 => "10111001",
 7812 => "01010101",
 7813 => "11110011",
 7814 => "10011001",
 7815 => "00001100",
 7816 => "01110010",
 7817 => "10010010",
 7818 => "00100100",
 7819 => "11100010",
 7820 => "01000110",
 7821 => "00110100",
 7822 => "11000001",
 7823 => "01111100",
 7824 => "10000101",
 7825 => "10000000",
 7826 => "11010001",
 7827 => "10110010",
 7828 => "10101000",
 7829 => "11100111",
 7830 => "11011010",
 7831 => "10011001",
 7832 => "00001011",
 7833 => "00100011",
 7834 => "10000111",
 7835 => "01001101",
 7836 => "11000101",
 7837 => "10101110",
 7838 => "00011111",
 7839 => "01010011",
 7840 => "00100011",
 7841 => "10111111",
 7842 => "11010110",
 7843 => "10111000",
 7844 => "10000000",
 7845 => "10000010",
 7846 => "01101100",
 7847 => "00111010",
 7848 => "01100010",
 7849 => "10100111",
 7850 => "10111110",
 7851 => "01110111",
 7852 => "10101010",
 7853 => "01100010",
 7854 => "00000011",
 7855 => "00111011",
 7856 => "00011001",
 7857 => "00101101",
 7858 => "11110000",
 7859 => "01110011",
 7860 => "00001111",
 7861 => "10111100",
 7862 => "11000000",
 7863 => "10010110",
 7864 => "10110100",
 7865 => "10101110",
 7866 => "01110011",
 7867 => "10100101",
 7868 => "11011110",
 7869 => "00101110",
 7870 => "11010100",
 7871 => "10100111",
 7872 => "01011111",
 7873 => "11100000",
 7874 => "01110010",
 7875 => "00111000",
 7876 => "10110000",
 7877 => "00000101",
 7878 => "00011000",
 7879 => "00111111",
 7880 => "10011011",
 7881 => "01110000",
 7882 => "10000110",
 7883 => "11010010",
 7884 => "00100001",
 7885 => "00000100",
 7886 => "01101011",
 7887 => "11100001",
 7888 => "11100001",
 7889 => "00010111",
 7890 => "01111010",
 7891 => "10001111",
 7892 => "11101001",
 7893 => "11001100",
 7894 => "01000110",
 7895 => "01011010",
 7896 => "01101110",
 7897 => "00010100",
 7898 => "11001010",
 7899 => "11011101",
 7900 => "10011000",
 7901 => "11100011",
 7902 => "01100110",
 7903 => "01100100",
 7904 => "00010101",
 7905 => "10100111",
 7906 => "01111110",
 7907 => "00010100",
 7908 => "11010100",
 7909 => "01000101",
 7910 => "11100010",
 7911 => "10111010",
 7912 => "01001100",
 7913 => "01100101",
 7914 => "00000110",
 7915 => "00001111",
 7916 => "00000100",
 7917 => "10101101",
 7918 => "10011101",
 7919 => "01111010",
 7920 => "01111011",
 7921 => "01101011",
 7922 => "11000010",
 7923 => "11001110",
 7924 => "00001101",
 7925 => "01110011",
 7926 => "10111010",
 7927 => "00111011",
 7928 => "11001010",
 7929 => "10101111",
 7930 => "00010010",
 7931 => "01100000",
 7932 => "01101111",
 7933 => "00110000",
 7934 => "11101011",
 7935 => "01001000",
 7936 => "00001100",
 7937 => "10011011",
 7938 => "10010011",
 7939 => "01111000",
 7940 => "11001010",
 7941 => "11011100",
 7942 => "10111111",
 7943 => "11000111",
 7944 => "00101100",
 7945 => "01000011",
 7946 => "11001001",
 7947 => "01110000",
 7948 => "11110111",
 7949 => "00101110",
 7950 => "11011110",
 7951 => "11010000",
 7952 => "00100111",
 7953 => "00001001",
 7954 => "00110000",
 7955 => "11111011",
 7956 => "10111010",
 7957 => "11111111",
 7958 => "00100001",
 7959 => "00001001",
 7960 => "10101110",
 7961 => "01100101",
 7962 => "10111011",
 7963 => "10010111",
 7964 => "11010010",
 7965 => "00011000",
 7966 => "10000101",
 7967 => "00110001",
 7968 => "01110011",
 7969 => "10101110",
 7970 => "11000000",
 7971 => "01010100",
 7972 => "11010001",
 7973 => "00011000",
 7974 => "01101011",
 7975 => "00101110",
 7976 => "00010101",
 7977 => "11011110",
 7978 => "11010110",
 7979 => "11111000",
 7980 => "01110101",
 7981 => "00111101",
 7982 => "01100010",
 7983 => "11110000",
 7984 => "10111101",
 7985 => "11100011",
 7986 => "00110100",
 7987 => "00000101",
 7988 => "10111110",
 7989 => "10101001",
 7990 => "10000011",
 7991 => "00101010",
 7992 => "10010101",
 7993 => "00110010",
 7994 => "01101000",
 7995 => "00100100",
 7996 => "10110110",
 7997 => "00100100",
 7998 => "10111100",
 7999 => "01010011",
 8000 => "11011001",
 8001 => "11101111",
 8002 => "01010011",
 8003 => "00010010",
 8004 => "00111111",
 8005 => "11010110",
 8006 => "00001111",
 8007 => "11000101",
 8008 => "00110001",
 8009 => "00100101",
 8010 => "00000010",
 8011 => "00110010",
 8012 => "01110111",
 8013 => "11000010",
 8014 => "11000100",
 8015 => "11111110",
 8016 => "00000011",
 8017 => "10101101",
 8018 => "00100000",
 8019 => "00010001",
 8020 => "11010000",
 8021 => "01011111",
 8022 => "10001100",
 8023 => "11001100",
 8024 => "01000010",
 8025 => "01111100",
 8026 => "01110000",
 8027 => "10010110",
 8028 => "00000000",
 8029 => "11110010",
 8030 => "11100101",
 8031 => "11001001",
 8032 => "11100010",
 8033 => "01100000",
 8034 => "01110111",
 8035 => "00100100",
 8036 => "11101001",
 8037 => "00110100",
 8038 => "11110010",
 8039 => "00110001",
 8040 => "10101101",
 8041 => "00101001",
 8042 => "00110001",
 8043 => "11110111",
 8044 => "11111101",
 8045 => "00001000",
 8046 => "01110011",
 8047 => "10011010",
 8048 => "10000011",
 8049 => "01001110",
 8050 => "00100101",
 8051 => "11001001",
 8052 => "11111001",
 8053 => "11011110",
 8054 => "10001100",
 8055 => "10110111",
 8056 => "11000111",
 8057 => "11100011",
 8058 => "11010010",
 8059 => "01111100",
 8060 => "01100011",
 8061 => "00100011",
 8062 => "01100001",
 8063 => "00111011",
 8064 => "10011100",
 8065 => "10001010",
 8066 => "00101011",
 8067 => "01100000",
 8068 => "10011100",
 8069 => "00100100",
 8070 => "00110100",
 8071 => "01101001",
 8072 => "10110000",
 8073 => "00111100",
 8074 => "01111100",
 8075 => "11100100",
 8076 => "11111001",
 8077 => "00101111",
 8078 => "11101101",
 8079 => "10101010",
 8080 => "00001110",
 8081 => "01110100",
 8082 => "11011100",
 8083 => "00011001",
 8084 => "10010010",
 8085 => "00001010",
 8086 => "00010001",
 8087 => "01011111",
 8088 => "00010100",
 8089 => "11000000",
 8090 => "01111100",
 8091 => "00111001",
 8092 => "00010101",
 8093 => "00110001",
 8094 => "10000111",
 8095 => "01010110",
 8096 => "00011110",
 8097 => "00100110",
 8098 => "01000101",
 8099 => "01000101",
 8100 => "00101100",
 8101 => "11010000",
 8102 => "00100100",
 8103 => "00101011",
 8104 => "00111100",
 8105 => "10001101",
 8106 => "10010101",
 8107 => "01110001",
 8108 => "01111111",
 8109 => "11101000",
 8110 => "01011001",
 8111 => "00111101",
 8112 => "00010101",
 8113 => "01110100",
 8114 => "10001010",
 8115 => "10111011",
 8116 => "00000100",
 8117 => "11111101",
 8118 => "01000101",
 8119 => "11011100",
 8120 => "00101100",
 8121 => "00111100",
 8122 => "00011110",
 8123 => "01101010",
 8124 => "01010111",
 8125 => "00110101",
 8126 => "01101011",
 8127 => "01110100",
 8128 => "11011101",
 8129 => "01101111",
 8130 => "10000101",
 8131 => "00011001",
 8132 => "01111111",
 8133 => "10001000",
 8134 => "01011111",
 8135 => "11110111",
 8136 => "01011011",
 8137 => "11000010",
 8138 => "10110111",
 8139 => "01111101",
 8140 => "00000001",
 8141 => "01010110",
 8142 => "01011011",
 8143 => "01110001",
 8144 => "00011000",
 8145 => "01001011",
 8146 => "11101001",
 8147 => "00101101",
 8148 => "00111011",
 8149 => "11001110",
 8150 => "01101001",
 8151 => "11001000",
 8152 => "10101101",
 8153 => "00111011",
 8154 => "11010000",
 8155 => "00000100",
 8156 => "01010001",
 8157 => "00110000",
 8158 => "00111100",
 8159 => "11011101",
 8160 => "10001001",
 8161 => "11011010",
 8162 => "01011100",
 8163 => "01010010",
 8164 => "11001101",
 8165 => "01011000",
 8166 => "01011110",
 8167 => "00010001",
 8168 => "00001100",
 8169 => "10011111",
 8170 => "00100100",
 8171 => "10011100",
 8172 => "00101010",
 8173 => "00001111",
 8174 => "01001000",
 8175 => "00011011",
 8176 => "01000101",
 8177 => "00000001",
 8178 => "10110001",
 8179 => "01000001",
 8180 => "11011101",
 8181 => "01100101",
 8182 => "11011000",
 8183 => "10001111",
 8184 => "11011010",
 8185 => "00001110",
 8186 => "11100110",
 8187 => "01011110",
 8188 => "11011111",
 8189 => "01000101",
 8190 => "01000001",
 8191 => "11010101",
 8192 => "11001101",
 8193 => "00110110",
 8194 => "10000111",
 8195 => "01100100",
 8196 => "00111001",
 8197 => "10001111",
 8198 => "11001001",
 8199 => "01001101",
 8200 => "10100111",
 8201 => "01000100",
 8202 => "10001000",
 8203 => "00001110",
 8204 => "10101111",
 8205 => "01011001",
 8206 => "01101010",
 8207 => "01001010",
 8208 => "01111101",
 8209 => "11111010",
 8210 => "01100010",
 8211 => "00000000",
 8212 => "10011111",
 8213 => "11011111",
 8214 => "11100011",
 8215 => "11101101",
 8216 => "01111100",
 8217 => "10100000",
 8218 => "11000101",
 8219 => "11101011",
 8220 => "10101111",
 8221 => "00000010",
 8222 => "01001000",
 8223 => "00000001",
 8224 => "11001101",
 8225 => "10000011",
 8226 => "01111011",
 8227 => "01100111",
 8228 => "11110001",
 8229 => "10101000",
 8230 => "10100111",
 8231 => "00001110",
 8232 => "10011111",
 8233 => "00100010",
 8234 => "10000111",
 8235 => "11111111",
 8236 => "00101100",
 8237 => "00110101",
 8238 => "00010111",
 8239 => "00111010",
 8240 => "01110011",
 8241 => "00101111",
 8242 => "00000100",
 8243 => "01011001",
 8244 => "00110101",
 8245 => "00000011",
 8246 => "11010000",
 8247 => "00001101",
 8248 => "00010100",
 8249 => "10101111",
 8250 => "11100010",
 8251 => "11000011",
 8252 => "00110010",
 8253 => "10010010",
 8254 => "01110011",
 8255 => "11111001",
 8256 => "00100110",
 8257 => "11011011",
 8258 => "10110001",
 8259 => "11110000",
 8260 => "01010001",
 8261 => "10110100",
 8262 => "01010011",
 8263 => "01011001",
 8264 => "10000111",
 8265 => "11000000",
 8266 => "10001111",
 8267 => "00000001",
 8268 => "10101111",
 8269 => "10000000",
 8270 => "00100000",
 8271 => "00010000",
 8272 => "11100000",
 8273 => "11101011",
 8274 => "11101010",
 8275 => "10011010",
 8276 => "11010001",
 8277 => "11110111",
 8278 => "00010000",
 8279 => "01110000",
 8280 => "10100111",
 8281 => "01110111",
 8282 => "10100010",
 8283 => "10011100",
 8284 => "01101101",
 8285 => "11010010",
 8286 => "01000011",
 8287 => "11101011",
 8288 => "11001000",
 8289 => "01100001",
 8290 => "00001000",
 8291 => "10110010",
 8292 => "11001111",
 8293 => "01001010",
 8294 => "10101111",
 8295 => "10000100",
 8296 => "10010111",
 8297 => "00111100",
 8298 => "01100001",
 8299 => "00100000",
 8300 => "11110101",
 8301 => "00110101",
 8302 => "10111100",
 8303 => "10110000",
 8304 => "01001011",
 8305 => "11101110",
 8306 => "11101101",
 8307 => "10001000",
 8308 => "00110000",
 8309 => "11101011",
 8310 => "11000011",
 8311 => "00001001",
 8312 => "10011011",
 8313 => "00101110",
 8314 => "01111000",
 8315 => "01000110",
 8316 => "10011001",
 8317 => "11101010",
 8318 => "00000101",
 8319 => "11100111",
 8320 => "11000110",
 8321 => "01110111",
 8322 => "00001100",
 8323 => "01000011",
 8324 => "01001100",
 8325 => "00010010",
 8326 => "11001101",
 8327 => "11110100",
 8328 => "01001011",
 8329 => "10010101",
 8330 => "01011110",
 8331 => "10011010",
 8332 => "00011010",
 8333 => "11010010",
 8334 => "00010100",
 8335 => "11101010",
 8336 => "01001000",
 8337 => "01010010",
 8338 => "10011101",
 8339 => "11101000",
 8340 => "11000010",
 8341 => "00011000",
 8342 => "10101010",
 8343 => "00101111",
 8344 => "10000000",
 8345 => "00101000",
 8346 => "10011010",
 8347 => "00011110",
 8348 => "01011100",
 8349 => "00001011",
 8350 => "01110001",
 8351 => "01100111",
 8352 => "10110011",
 8353 => "10011001",
 8354 => "11100010",
 8355 => "10110101",
 8356 => "00111110",
 8357 => "01011001",
 8358 => "10110010",
 8359 => "10111010",
 8360 => "10001010",
 8361 => "11010110",
 8362 => "11010010",
 8363 => "10011101",
 8364 => "10100110",
 8365 => "00010001",
 8366 => "01100010",
 8367 => "11111101",
 8368 => "10011111",
 8369 => "10100100",
 8370 => "01010100",
 8371 => "10010001",
 8372 => "00100010",
 8373 => "10110001",
 8374 => "11101100",
 8375 => "11001010",
 8376 => "00000011",
 8377 => "00000111",
 8378 => "10000011",
 8379 => "01111100",
 8380 => "01111110",
 8381 => "01110001",
 8382 => "01111001",
 8383 => "10101010",
 8384 => "01001010",
 8385 => "11100001",
 8386 => "11010111",
 8387 => "11011111",
 8388 => "01100110",
 8389 => "11000011",
 8390 => "01111110",
 8391 => "11100011",
 8392 => "10001010",
 8393 => "11100000",
 8394 => "01110111",
 8395 => "11001100",
 8396 => "11011111",
 8397 => "01000011",
 8398 => "10011100",
 8399 => "01001100",
 8400 => "01000011",
 8401 => "00011011",
 8402 => "00100001",
 8403 => "01110111",
 8404 => "00001110",
 8405 => "10000101",
 8406 => "00111111",
 8407 => "01101000",
 8408 => "01010101",
 8409 => "00101011",
 8410 => "10100100",
 8411 => "11010000",
 8412 => "11110001",
 8413 => "00110100",
 8414 => "01101100",
 8415 => "00111000",
 8416 => "11011010",
 8417 => "00010101",
 8418 => "10011110",
 8419 => "10100101",
 8420 => "10101101",
 8421 => "11110101",
 8422 => "00000001",
 8423 => "00101110",
 8424 => "00011110",
 8425 => "01101111",
 8426 => "10010000",
 8427 => "00110000",
 8428 => "11110000",
 8429 => "10101100",
 8430 => "00010110",
 8431 => "11000100",
 8432 => "10100011",
 8433 => "00011010",
 8434 => "11011110",
 8435 => "01001001",
 8436 => "01011011",
 8437 => "11000111",
 8438 => "01111000",
 8439 => "11001011",
 8440 => "11000110",
 8441 => "11110010",
 8442 => "11101001",
 8443 => "10111100",
 8444 => "11011001",
 8445 => "00001101",
 8446 => "11110000",
 8447 => "00001010",
 8448 => "11000110",
 8449 => "11000000",
 8450 => "01110101",
 8451 => "00011101",
 8452 => "11010110",
 8453 => "00011000",
 8454 => "01001111",
 8455 => "00101010",
 8456 => "10101000",
 8457 => "10001100",
 8458 => "01101010",
 8459 => "10000000",
 8460 => "00110111",
 8461 => "10000100",
 8462 => "00010000",
 8463 => "11010100",
 8464 => "10111000",
 8465 => "10011101",
 8466 => "10011110",
 8467 => "00111001",
 8468 => "10111010",
 8469 => "11001001",
 8470 => "00110111",
 8471 => "11000010",
 8472 => "01100110",
 8473 => "11001000",
 8474 => "10001011",
 8475 => "00110010",
 8476 => "00110100",
 8477 => "11011110",
 8478 => "11010010",
 8479 => "00011110",
 8480 => "10011100",
 8481 => "01010001",
 8482 => "01111111",
 8483 => "10000110",
 8484 => "10010000",
 8485 => "01001001",
 8486 => "01110011",
 8487 => "00110011",
 8488 => "01101011",
 8489 => "01010110",
 8490 => "10001111",
 8491 => "00010110",
 8492 => "00000111",
 8493 => "01000011",
 8494 => "11001110",
 8495 => "01000100",
 8496 => "10100101",
 8497 => "11011100",
 8498 => "01100100",
 8499 => "00000010",
 8500 => "01001100",
 8501 => "11001001",
 8502 => "01011001",
 8503 => "01100000",
 8504 => "01110110",
 8505 => "10010110",
 8506 => "11011101",
 8507 => "11000011",
 8508 => "00011111",
 8509 => "11010010",
 8510 => "11100000",
 8511 => "01100110",
 8512 => "11000100",
 8513 => "10101100",
 8514 => "01101011",
 8515 => "11010100",
 8516 => "01000011",
 8517 => "11001000",
 8518 => "00100010",
 8519 => "10001110",
 8520 => "10100000",
 8521 => "10000110",
 8522 => "11110101",
 8523 => "11011100",
 8524 => "01000010",
 8525 => "10001101",
 8526 => "10100111",
 8527 => "01111110",
 8528 => "00010111",
 8529 => "00011100",
 8530 => "11110111",
 8531 => "00011010",
 8532 => "10000000",
 8533 => "00110110",
 8534 => "00010100",
 8535 => "10000101",
 8536 => "10111000",
 8537 => "10111111",
 8538 => "01110101",
 8539 => "00101010",
 8540 => "10011011",
 8541 => "00100001",
 8542 => "10010011",
 8543 => "00101110",
 8544 => "01101100",
 8545 => "11111101",
 8546 => "10001001",
 8547 => "00100101",
 8548 => "11101000",
 8549 => "00100011",
 8550 => "00101101",
 8551 => "11110000",
 8552 => "10010000",
 8553 => "10001010",
 8554 => "10101011",
 8555 => "01111000",
 8556 => "00110011",
 8557 => "10101001",
 8558 => "11110011",
 8559 => "01100001",
 8560 => "01011101",
 8561 => "11000000",
 8562 => "10101000",
 8563 => "00010000",
 8564 => "10100110",
 8565 => "00010010",
 8566 => "10101000",
 8567 => "00011010",
 8568 => "01011001",
 8569 => "11010110",
 8570 => "00101011",
 8571 => "11011110",
 8572 => "11000110",
 8573 => "01110110",
 8574 => "10100000",
 8575 => "01110110",
 8576 => "10111011",
 8577 => "10011100",
 8578 => "11010101",
 8579 => "10100010",
 8580 => "11110101",
 8581 => "10010001",
 8582 => "01010000",
 8583 => "11000000",
 8584 => "10101001",
 8585 => "01010000",
 8586 => "01010100",
 8587 => "11110011",
 8588 => "10100101",
 8589 => "10000110",
 8590 => "10001111",
 8591 => "10010100",
 8592 => "00010001",
 8593 => "00101101",
 8594 => "10100111",
 8595 => "00111000",
 8596 => "01010011",
 8597 => "11111110",
 8598 => "01100100",
 8599 => "01010100",
 8600 => "00100101",
 8601 => "01011101",
 8602 => "10101110",
 8603 => "10001110",
 8604 => "10001001",
 8605 => "11111011",
 8606 => "10100000",
 8607 => "01101110",
 8608 => "10010000",
 8609 => "11010111",
 8610 => "11110111",
 8611 => "10001110",
 8612 => "01011111",
 8613 => "10011001",
 8614 => "00101011",
 8615 => "00111101",
 8616 => "11000101",
 8617 => "00101011",
 8618 => "10111000",
 8619 => "10010000",
 8620 => "01001101",
 8621 => "10011111",
 8622 => "00011100",
 8623 => "00000010",
 8624 => "01000111",
 8625 => "11100101",
 8626 => "01011100",
 8627 => "10000000",
 8628 => "10100101",
 8629 => "11000010",
 8630 => "01111100",
 8631 => "01110100",
 8632 => "10000101",
 8633 => "11101101",
 8634 => "11110000",
 8635 => "11000001",
 8636 => "01100100",
 8637 => "00010010",
 8638 => "00101010",
 8639 => "10110010",
 8640 => "00111000",
 8641 => "11001100",
 8642 => "00101101",
 8643 => "11111111",
 8644 => "00001010",
 8645 => "01100100",
 8646 => "10011101",
 8647 => "01010000",
 8648 => "10001010",
 8649 => "10001100",
 8650 => "11100111",
 8651 => "11001000",
 8652 => "01100110",
 8653 => "11001010",
 8654 => "00110100",
 8655 => "11010000",
 8656 => "11111011",
 8657 => "01010011",
 8658 => "11101011",
 8659 => "01101101",
 8660 => "01011101",
 8661 => "00101000",
 8662 => "10110000",
 8663 => "11100111",
 8664 => "00000110",
 8665 => "11111000",
 8666 => "01010101",
 8667 => "10111001",
 8668 => "01001111",
 8669 => "00010010",
 8670 => "10100000",
 8671 => "10001111",
 8672 => "01100011",
 8673 => "11111101",
 8674 => "11000100",
 8675 => "10010101",
 8676 => "11100000",
 8677 => "10000101",
 8678 => "10101001",
 8679 => "01111000",
 8680 => "00110110",
 8681 => "00000101",
 8682 => "01010111",
 8683 => "00000111",
 8684 => "00100001",
 8685 => "11110111",
 8686 => "01000111",
 8687 => "00110101",
 8688 => "10111000",
 8689 => "11010101",
 8690 => "10100101",
 8691 => "10001110",
 8692 => "11001011",
 8693 => "10100011",
 8694 => "11111011",
 8695 => "11111100",
 8696 => "00101111",
 8697 => "00000000",
 8698 => "01000100",
 8699 => "11110011",
 8700 => "10000001",
 8701 => "00001010",
 8702 => "00010000",
 8703 => "10011100",
 8704 => "00000110",
 8705 => "10110011",
 8706 => "00100001",
 8707 => "01001101",
 8708 => "10011000",
 8709 => "11000100",
 8710 => "00011110",
 8711 => "10000011",
 8712 => "11001011",
 8713 => "11100101",
 8714 => "01011001",
 8715 => "01110000",
 8716 => "10011100",
 8717 => "11110000",
 8718 => "11101001",
 8719 => "00101000",
 8720 => "11011001",
 8721 => "10010000",
 8722 => "01011110",
 8723 => "01011101",
 8724 => "11010000",
 8725 => "01000000",
 8726 => "10011010",
 8727 => "01101100",
 8728 => "01110100",
 8729 => "10111111",
 8730 => "11100100",
 8731 => "11010100",
 8732 => "00111111",
 8733 => "00101001",
 8734 => "10110001",
 8735 => "01000111",
 8736 => "11000100",
 8737 => "11101001",
 8738 => "00101100",
 8739 => "00001011",
 8740 => "00000101",
 8741 => "01000111",
 8742 => "10100010",
 8743 => "10101101",
 8744 => "01111101",
 8745 => "11000101",
 8746 => "10111000",
 8747 => "11100101",
 8748 => "00010000",
 8749 => "11000011",
 8750 => "01010001",
 8751 => "00010110",
 8752 => "10010100",
 8753 => "11110010",
 8754 => "00100110",
 8755 => "00010010",
 8756 => "11111001",
 8757 => "01001000",
 8758 => "11111110",
 8759 => "00000111",
 8760 => "00001110",
 8761 => "00101001",
 8762 => "01101010",
 8763 => "01001111",
 8764 => "01011011",
 8765 => "01000110",
 8766 => "00001001",
 8767 => "01111111",
 8768 => "00100010",
 8769 => "00111101",
 8770 => "01000110",
 8771 => "11011100",
 8772 => "01011011",
 8773 => "10111010",
 8774 => "10111110",
 8775 => "01100101",
 8776 => "00000001",
 8777 => "10100100",
 8778 => "01001101",
 8779 => "01000110",
 8780 => "01110110",
 8781 => "10011010",
 8782 => "00110001",
 8783 => "11111010",
 8784 => "00101110",
 8785 => "01001111",
 8786 => "10111110",
 8787 => "10000011",
 8788 => "11001010",
 8789 => "01110001",
 8790 => "10101111",
 8791 => "01011000",
 8792 => "00110100",
 8793 => "01001000",
 8794 => "01110010",
 8795 => "01101100",
 8796 => "01010010",
 8797 => "01100101",
 8798 => "01110000",
 8799 => "00101111",
 8800 => "10111100",
 8801 => "10101111",
 8802 => "01011010",
 8803 => "00001100",
 8804 => "11011011",
 8805 => "10001101",
 8806 => "11011010",
 8807 => "01010001",
 8808 => "01011101",
 8809 => "10110101",
 8810 => "11011011",
 8811 => "00010110",
 8812 => "10100010",
 8813 => "11000111",
 8814 => "11010101",
 8815 => "10011010",
 8816 => "00010000",
 8817 => "11111110",
 8818 => "01111010",
 8819 => "01010110",
 8820 => "00010001",
 8821 => "01100000",
 8822 => "11000101",
 8823 => "11001010",
 8824 => "10000100",
 8825 => "01110101",
 8826 => "01001001",
 8827 => "00000010",
 8828 => "01011111",
 8829 => "11100000",
 8830 => "11111000",
 8831 => "00101111",
 8832 => "00011111",
 8833 => "00101101",
 8834 => "00111001",
 8835 => "00100010",
 8836 => "11010111",
 8837 => "00000011",
 8838 => "01110011",
 8839 => "11101111",
 8840 => "10101010",
 8841 => "11011100",
 8842 => "01100000",
 8843 => "11100011",
 8844 => "11101001",
 8845 => "00110101",
 8846 => "01111111",
 8847 => "10010100",
 8848 => "10111101",
 8849 => "11010110",
 8850 => "01111101",
 8851 => "01110001",
 8852 => "00010001",
 8853 => "10010110",
 8854 => "10110010",
 8855 => "00111001",
 8856 => "00010100",
 8857 => "00000111",
 8858 => "11111000",
 8859 => "00001011",
 8860 => "01011110",
 8861 => "11011011",
 8862 => "11000011",
 8863 => "00010010",
 8864 => "10100111",
 8865 => "00100001",
 8866 => "10110110",
 8867 => "01111100",
 8868 => "10111110",
 8869 => "11110110",
 8870 => "01010001",
 8871 => "10110011",
 8872 => "00010101",
 8873 => "10101111",
 8874 => "01011101",
 8875 => "00011110",
 8876 => "00010100",
 8877 => "01011000",
 8878 => "00010110",
 8879 => "00111000",
 8880 => "00110001",
 8881 => "00101100",
 8882 => "11011111",
 8883 => "11000000",
 8884 => "00011001",
 8885 => "10100100",
 8886 => "01111001",
 8887 => "00011110",
 8888 => "01110110",
 8889 => "01101110",
 8890 => "10010110",
 8891 => "10101000",
 8892 => "01000010",
 8893 => "01110110",
 8894 => "00010011",
 8895 => "10011010",
 8896 => "00111010",
 8897 => "00101001",
 8898 => "01011001",
 8899 => "00001000",
 8900 => "00101000",
 8901 => "01011000",
 8902 => "11000110",
 8903 => "10000101",
 8904 => "11001101",
 8905 => "01001000",
 8906 => "01010010",
 8907 => "11110101",
 8908 => "01111100",
 8909 => "11100011",
 8910 => "11001010",
 8911 => "00001001",
 8912 => "01010000",
 8913 => "00001000",
 8914 => "01011001",
 8915 => "11001110",
 8916 => "00100001",
 8917 => "01110111",
 8918 => "00001000",
 8919 => "10011110",
 8920 => "11100100",
 8921 => "01110001",
 8922 => "11110001",
 8923 => "10010101",
 8924 => "10111110",
 8925 => "10001100",
 8926 => "01100000",
 8927 => "00001101",
 8928 => "00011011",
 8929 => "11010101",
 8930 => "11010111",
 8931 => "01111111",
 8932 => "11010011",
 8933 => "00100001",
 8934 => "00100100",
 8935 => "10010101",
 8936 => "10000000",
 8937 => "01111111",
 8938 => "11100101",
 8939 => "00000000",
 8940 => "10001010",
 8941 => "01011100",
 8942 => "01101000",
 8943 => "10110011",
 8944 => "01100000",
 8945 => "00011010",
 8946 => "00010011",
 8947 => "10011011",
 8948 => "10110010",
 8949 => "10111101",
 8950 => "11000101",
 8951 => "10110001",
 8952 => "11100111",
 8953 => "10100001",
 8954 => "00000000",
 8955 => "10101000",
 8956 => "01100111",
 8957 => "11001010",
 8958 => "11110001",
 8959 => "00010100",
 8960 => "10001111",
 8961 => "01100101",
 8962 => "11001101",
 8963 => "10001100",
 8964 => "10101110",
 8965 => "01110010",
 8966 => "01010101",
 8967 => "00111011",
 8968 => "01000010",
 8969 => "11100111",
 8970 => "01101000",
 8971 => "00010101",
 8972 => "11100101",
 8973 => "11111000",
 8974 => "01101010",
 8975 => "11011000",
 8976 => "11001010",
 8977 => "01000110",
 8978 => "10100110",
 8979 => "11101000",
 8980 => "00001101",
 8981 => "00110000",
 8982 => "01010000",
 8983 => "00001111",
 8984 => "11101000",
 8985 => "10001001",
 8986 => "10001101",
 8987 => "00011100",
 8988 => "00001111",
 8989 => "10110010",
 8990 => "10010110",
 8991 => "00001110",
 8992 => "01010000",
 8993 => "10001111",
 8994 => "11100001",
 8995 => "01100110",
 8996 => "00110111",
 8997 => "10110101",
 8998 => "01100000",
 8999 => "01000010",
 9000 => "01100110",
 9001 => "00111111",
 9002 => "11100100",
 9003 => "00110100",
 9004 => "10100100",
 9005 => "11101101",
 9006 => "10001000",
 9007 => "11011101",
 9008 => "11110010",
 9009 => "11111111",
 9010 => "01000011",
 9011 => "11111000",
 9012 => "11001110",
 9013 => "11101110",
 9014 => "00100011",
 9015 => "11100111",
 9016 => "10100110",
 9017 => "00001111",
 9018 => "10101000",
 9019 => "11001111",
 9020 => "10111100",
 9021 => "10100110",
 9022 => "00001101",
 9023 => "01101101",
 9024 => "10110001",
 9025 => "00001000",
 9026 => "01101001",
 9027 => "00011011",
 9028 => "10100100",
 9029 => "11100101",
 9030 => "00011000",
 9031 => "11110101",
 9032 => "10100011",
 9033 => "01101110",
 9034 => "10101001",
 9035 => "01010101",
 9036 => "01110010",
 9037 => "01001001",
 9038 => "10111010",
 9039 => "00111010",
 9040 => "11111110",
 9041 => "01010100",
 9042 => "00100001",
 9043 => "01110111",
 9044 => "10100010",
 9045 => "01111001",
 9046 => "10111010",
 9047 => "00100100",
 9048 => "01000000",
 9049 => "00110010",
 9050 => "11010001",
 9051 => "11011000",
 9052 => "11101111",
 9053 => "00110000",
 9054 => "01001101",
 9055 => "10001000",
 9056 => "10000000",
 9057 => "11111010",
 9058 => "01110111",
 9059 => "00101010",
 9060 => "10110110",
 9061 => "01010010",
 9062 => "10011000",
 9063 => "01001000",
 9064 => "01100100",
 9065 => "01111111",
 9066 => "11011010",
 9067 => "01001010",
 9068 => "10001111",
 9069 => "01100111",
 9070 => "00101010",
 9071 => "00110011",
 9072 => "01000111",
 9073 => "00100000",
 9074 => "11111010",
 9075 => "01010111",
 9076 => "01110110",
 9077 => "11100010",
 9078 => "11010011",
 9079 => "01011110",
 9080 => "10000000",
 9081 => "00001000",
 9082 => "10110100",
 9083 => "00111100",
 9084 => "10111100",
 9085 => "11100011",
 9086 => "01110110",
 9087 => "00100010",
 9088 => "01000000",
 9089 => "11001011",
 9090 => "10110111",
 9091 => "10011100",
 9092 => "00010101",
 9093 => "11010111",
 9094 => "01100010",
 9095 => "11110111",
 9096 => "00110101",
 9097 => "01110011",
 9098 => "10000111",
 9099 => "11110010",
 9100 => "10010111",
 9101 => "00110000",
 9102 => "10010001",
 9103 => "01101101",
 9104 => "01111101",
 9105 => "10011011",
 9106 => "11000010",
 9107 => "11111111",
 9108 => "10000110",
 9109 => "11100001",
 9110 => "01110000",
 9111 => "11111111",
 9112 => "11011011",
 9113 => "00101010",
 9114 => "11000000",
 9115 => "00111000",
 9116 => "01101111",
 9117 => "10000011",
 9118 => "00111011",
 9119 => "00100101",
 9120 => "01000011",
 9121 => "11000000",
 9122 => "00011101",
 9123 => "10001011",
 9124 => "11101010",
 9125 => "01010010",
 9126 => "01101000",
 9127 => "11000010",
 9128 => "00010000",
 9129 => "01111110",
 9130 => "11000110",
 9131 => "01010111",
 9132 => "01110101",
 9133 => "10011111",
 9134 => "00000100",
 9135 => "00100100",
 9136 => "01101001",
 9137 => "01001001",
 9138 => "10001000",
 9139 => "01000001",
 9140 => "10001111",
 9141 => "11011001",
 9142 => "10001101",
 9143 => "10010110",
 9144 => "10111011",
 9145 => "00110111",
 9146 => "10011110",
 9147 => "11001110",
 9148 => "10111000",
 9149 => "10111100",
 9150 => "01001101",
 9151 => "01100101",
 9152 => "01001000",
 9153 => "11101001",
 9154 => "10000010",
 9155 => "11000111",
 9156 => "01100111",
 9157 => "11000101",
 9158 => "01101011",
 9159 => "00010101",
 9160 => "11100010",
 9161 => "01101001",
 9162 => "01101000",
 9163 => "11111110",
 9164 => "10110101",
 9165 => "11100010",
 9166 => "00110101",
 9167 => "10000000",
 9168 => "10000100",
 9169 => "10111110",
 9170 => "01100000",
 9171 => "11110111",
 9172 => "10001111",
 9173 => "00110010",
 9174 => "01001110",
 9175 => "10100001",
 9176 => "11000111",
 9177 => "10011010",
 9178 => "10010011",
 9179 => "11011100",
 9180 => "00000010",
 9181 => "11111111",
 9182 => "01001000",
 9183 => "01001000",
 9184 => "01011110",
 9185 => "10100101",
 9186 => "11100001",
 9187 => "01100000",
 9188 => "01111111",
 9189 => "00100101",
 9190 => "00111010",
 9191 => "10001111",
 9192 => "10011110",
 9193 => "01100111",
 9194 => "00000000",
 9195 => "11011110",
 9196 => "11110010",
 9197 => "10010011",
 9198 => "01101100",
 9199 => "11000011",
 9200 => "00101101",
 9201 => "01111100",
 9202 => "10110011",
 9203 => "01011101",
 9204 => "11010000",
 9205 => "11010010",
 9206 => "00011001",
 9207 => "01101111",
 9208 => "00011000",
 9209 => "10111110",
 9210 => "00110000",
 9211 => "11000001",
 9212 => "10010001",
 9213 => "00001011",
 9214 => "10111110",
 9215 => "00101111",
 9216 => "10000000",
 9217 => "11000011",
 9218 => "11111101",
 9219 => "00100001",
 9220 => "10001100",
 9221 => "00100111",
 9222 => "10101001",
 9223 => "00100011",
 9224 => "10100001",
 9225 => "00101111",
 9226 => "00011010",
 9227 => "01110001",
 9228 => "11011011",
 9229 => "01100010",
 9230 => "10101101",
 9231 => "10011100",
 9232 => "00110101",
 9233 => "01000011",
 9234 => "11111110",
 9235 => "01000010",
 9236 => "00110011",
 9237 => "00001110",
 9238 => "11110011",
 9239 => "00001111",
 9240 => "11000110",
 9241 => "11011100",
 9242 => "01111100",
 9243 => "11010000",
 9244 => "00110000",
 9245 => "00000111",
 9246 => "01000111",
 9247 => "10011111",
 9248 => "10011000",
 9249 => "01001101",
 9250 => "11010000",
 9251 => "10101010",
 9252 => "01000111",
 9253 => "10100101",
 9254 => "11111111",
 9255 => "11010101",
 9256 => "01111100",
 9257 => "10110000",
 9258 => "11010100",
 9259 => "11111001",
 9260 => "01111010",
 9261 => "11001101",
 9262 => "00111110",
 9263 => "01010111",
 9264 => "00110011",
 9265 => "00001111",
 9266 => "00001110",
 9267 => "00100111",
 9268 => "01110101",
 9269 => "01111011",
 9270 => "00101011",
 9271 => "00111010",
 9272 => "11101101",
 9273 => "01011100",
 9274 => "10010010",
 9275 => "11100000",
 9276 => "10110001",
 9277 => "00101100",
 9278 => "10011110",
 9279 => "00010100",
 9280 => "11000100",
 9281 => "01111010",
 9282 => "11111110",
 9283 => "10000110",
 9284 => "00111010",
 9285 => "10011110",
 9286 => "00100110",
 9287 => "01110010",
 9288 => "00111010",
 9289 => "11111011",
 9290 => "11111011",
 9291 => "00000111",
 9292 => "10110101",
 9293 => "01011110",
 9294 => "00001100",
 9295 => "11011100",
 9296 => "01100101",
 9297 => "00001010",
 9298 => "01110111",
 9299 => "11000000",
 9300 => "11110100",
 9301 => "11001101",
 9302 => "10000101",
 9303 => "00000000",
 9304 => "00100011",
 9305 => "10101111",
 9306 => "01111010",
 9307 => "01010010",
 9308 => "00000111",
 9309 => "10100100",
 9310 => "01111100",
 9311 => "11001100",
 9312 => "00000111",
 9313 => "11001100",
 9314 => "11010011",
 9315 => "00101111",
 9316 => "11100001",
 9317 => "10010001",
 9318 => "00110111",
 9319 => "00001010",
 9320 => "10111100",
 9321 => "00101011",
 9322 => "10011000",
 9323 => "10111100",
 9324 => "10101011",
 9325 => "00001001",
 9326 => "11110001",
 9327 => "11100101",
 9328 => "11000111",
 9329 => "00101000",
 9330 => "00011000",
 9331 => "00010011",
 9332 => "01011010",
 9333 => "11010110",
 9334 => "10100010",
 9335 => "10111001",
 9336 => "10010111",
 9337 => "11000111",
 9338 => "11001100",
 9339 => "01111111",
 9340 => "11011011",
 9341 => "11001011",
 9342 => "11110101",
 9343 => "10101000",
 9344 => "01010000",
 9345 => "00111110",
 9346 => "10110010",
 9347 => "11101001",
 9348 => "00000010",
 9349 => "00010000",
 9350 => "11101100",
 9351 => "11111000",
 9352 => "10001101",
 9353 => "10110001",
 9354 => "01111011",
 9355 => "00011101",
 9356 => "10111011",
 9357 => "10101000",
 9358 => "10010001",
 9359 => "00010111",
 9360 => "11110001",
 9361 => "11010100",
 9362 => "11101111",
 9363 => "10100110",
 9364 => "10011110",
 9365 => "11001100",
 9366 => "00010110",
 9367 => "10110110",
 9368 => "01100100",
 9369 => "10100010",
 9370 => "01001110",
 9371 => "11101001",
 9372 => "01000111",
 9373 => "00000101",
 9374 => "00000010",
 9375 => "11010111",
 9376 => "01100100",
 9377 => "11100011",
 9378 => "10001001",
 9379 => "01011000",
 9380 => "11111101",
 9381 => "11010011",
 9382 => "11000110",
 9383 => "01111000",
 9384 => "11001111",
 9385 => "10001001",
 9386 => "11110000",
 9387 => "10001100",
 9388 => "01110011",
 9389 => "11010111",
 9390 => "01010111",
 9391 => "10111010",
 9392 => "01000110",
 9393 => "10000000",
 9394 => "00111010",
 9395 => "11001001",
 9396 => "00010010",
 9397 => "10011011",
 9398 => "00100111",
 9399 => "11111111",
 9400 => "00001010",
 9401 => "01000110",
 9402 => "10001110",
 9403 => "11010010",
 9404 => "11111001",
 9405 => "10101101",
 9406 => "11111011",
 9407 => "11001000",
 9408 => "01010100",
 9409 => "01111001",
 9410 => "00010011",
 9411 => "00001100",
 9412 => "10011010",
 9413 => "00010100",
 9414 => "00010110",
 9415 => "00000110",
 9416 => "01110011",
 9417 => "01101110",
 9418 => "01011111",
 9419 => "11010001",
 9420 => "01000000",
 9421 => "10100011",
 9422 => "10100010",
 9423 => "10101110",
 9424 => "11000011",
 9425 => "10011010",
 9426 => "11011101",
 9427 => "00110110",
 9428 => "11111010",
 9429 => "00011101",
 9430 => "10000000",
 9431 => "11110010",
 9432 => "01011001",
 9433 => "10100101",
 9434 => "01100100",
 9435 => "01111101",
 9436 => "11001001",
 9437 => "10001110",
 9438 => "11101001",
 9439 => "01000110",
 9440 => "11101111",
 9441 => "10001010",
 9442 => "11001110",
 9443 => "00100100",
 9444 => "00001000",
 9445 => "00100101",
 9446 => "10111111",
 9447 => "11110000",
 9448 => "00010001",
 9449 => "10100010",
 9450 => "10100110",
 9451 => "00010000",
 9452 => "00011000",
 9453 => "10011111",
 9454 => "10001011",
 9455 => "00001100",
 9456 => "11110011",
 9457 => "10011001",
 9458 => "10001110",
 9459 => "00010010",
 9460 => "00100111",
 9461 => "00100100",
 9462 => "00010111",
 9463 => "10100011",
 9464 => "10000000",
 9465 => "00001011",
 9466 => "11111010",
 9467 => "01101111",
 9468 => "10111101",
 9469 => "01011111",
 9470 => "10111010",
 9471 => "00111001",
 9472 => "10001011",
 9473 => "00001000",
 9474 => "10001001",
 9475 => "00110001",
 9476 => "11111111",
 9477 => "01011001",
 9478 => "01100101",
 9479 => "11101101",
 9480 => "00110100",
 9481 => "00011000",
 9482 => "10111110",
 9483 => "00000110",
 9484 => "10101011",
 9485 => "11110000",
 9486 => "01011011",
 9487 => "11011111",
 9488 => "00010111",
 9489 => "11111101",
 9490 => "11001011",
 9491 => "01010111",
 9492 => "10001100",
 9493 => "11000110",
 9494 => "01000111",
 9495 => "00000011",
 9496 => "01101010",
 9497 => "11011101",
 9498 => "11001000",
 9499 => "11001101",
 9500 => "01001010",
 9501 => "10000001",
 9502 => "10110000",
 9503 => "01110001",
 9504 => "01000100",
 9505 => "01111011",
 9506 => "10011010",
 9507 => "11100000",
 9508 => "10000111",
 9509 => "01010101",
 9510 => "00011100",
 9511 => "01111110",
 9512 => "01000110",
 9513 => "11111110",
 9514 => "11001101",
 9515 => "01010001",
 9516 => "11101010",
 9517 => "00110011",
 9518 => "01101010",
 9519 => "01010010",
 9520 => "10100101",
 9521 => "01001100",
 9522 => "00111011",
 9523 => "01000101",
 9524 => "01010101",
 9525 => "01000111",
 9526 => "10100100",
 9527 => "01000100",
 9528 => "11010000",
 9529 => "00101010",
 9530 => "00100000",
 9531 => "01100100",
 9532 => "10110011",
 9533 => "10100010",
 9534 => "01000110",
 9535 => "01001010",
 9536 => "10011011",
 9537 => "01000110",
 9538 => "11000100",
 9539 => "00110110",
 9540 => "11101001",
 9541 => "01100001",
 9542 => "10110010",
 9543 => "11110000",
 9544 => "11111010",
 9545 => "00110100",
 9546 => "10110110",
 9547 => "01111011",
 9548 => "11001111",
 9549 => "01001100",
 9550 => "00100110",
 9551 => "10000111",
 9552 => "01001000",
 9553 => "11111110",
 9554 => "01010100",
 9555 => "01110011",
 9556 => "01101101",
 9557 => "00110100",
 9558 => "10100101",
 9559 => "00000111",
 9560 => "10111110",
 9561 => "11011000",
 9562 => "00101011",
 9563 => "11001000",
 9564 => "10010110",
 9565 => "00100001",
 9566 => "00110100",
 9567 => "11011000",
 9568 => "00000010",
 9569 => "10011011",
 9570 => "10110010",
 9571 => "01011111",
 9572 => "10101000",
 9573 => "11011111",
 9574 => "10000011",
 9575 => "11011111",
 9576 => "01000011",
 9577 => "10000000",
 9578 => "01000000",
 9579 => "11100111",
 9580 => "11000001",
 9581 => "10001011",
 9582 => "11101011",
 9583 => "11011100",
 9584 => "10001011",
 9585 => "11001110",
 9586 => "11001110",
 9587 => "00001001",
 9588 => "10001110",
 9589 => "11100010",
 9590 => "00110011",
 9591 => "01010001",
 9592 => "10000100",
 9593 => "10010000",
 9594 => "11101011",
 9595 => "01100101",
 9596 => "00011110",
 9597 => "10110110",
 9598 => "00111011",
 9599 => "10100100",
 9600 => "01111101",
 9601 => "11110110",
 9602 => "00010111",
 9603 => "10111010",
 9604 => "10010101",
 9605 => "11001100",
 9606 => "01111101",
 9607 => "10010100",
 9608 => "01011110",
 9609 => "00001110",
 9610 => "11100111",
 9611 => "00001110",
 9612 => "00010011",
 9613 => "10110111",
 9614 => "11101101",
 9615 => "01101010",
 9616 => "11011111",
 9617 => "01010010",
 9618 => "11010000",
 9619 => "01111011",
 9620 => "01010110",
 9621 => "10010101",
 9622 => "01110010",
 9623 => "00110111",
 9624 => "10101010",
 9625 => "01001110",
 9626 => "11111010",
 9627 => "00101010",
 9628 => "01010010",
 9629 => "10000110",
 9630 => "11111011",
 9631 => "10011111",
 9632 => "00000111",
 9633 => "11000010",
 9634 => "10100001",
 9635 => "01010110",
 9636 => "01101100",
 9637 => "11001010",
 9638 => "11100000",
 9639 => "00001001",
 9640 => "11110111",
 9641 => "11101101",
 9642 => "00100111",
 9643 => "01100101",
 9644 => "00100010",
 9645 => "11100011",
 9646 => "11101111",
 9647 => "00001100",
 9648 => "11001010",
 9649 => "00010010",
 9650 => "11101100",
 9651 => "00111101",
 9652 => "00111011",
 9653 => "00110101",
 9654 => "11000111",
 9655 => "11110000",
 9656 => "01110010",
 9657 => "00000100",
 9658 => "10011000",
 9659 => "00000110",
 9660 => "11110111",
 9661 => "00100001",
 9662 => "10101000",
 9663 => "10100111",
 9664 => "00111111",
 9665 => "00011100",
 9666 => "11000110",
 9667 => "01011001",
 9668 => "00001001",
 9669 => "00101011",
 9670 => "00010000",
 9671 => "10111001",
 9672 => "00110011",
 9673 => "00100101",
 9674 => "01101010",
 9675 => "00001101",
 9676 => "01111010",
 9677 => "01010001",
 9678 => "00101100",
 9679 => "01111100",
 9680 => "01101101",
 9681 => "01010001",
 9682 => "00100101",
 9683 => "10011010",
 9684 => "00010010",
 9685 => "00000000",
 9686 => "11111111",
 9687 => "11101000",
 9688 => "00101100",
 9689 => "00110010",
 9690 => "10110100",
 9691 => "01010111",
 9692 => "01010000",
 9693 => "00010010",
 9694 => "11000000",
 9695 => "00110110",
 9696 => "10011001",
 9697 => "11010100",
 9698 => "10010110",
 9699 => "11000000",
 9700 => "01000000",
 9701 => "11101110",
 9702 => "00100100",
 9703 => "10011101",
 9704 => "01011001",
 9705 => "10011010",
 9706 => "00000100",
 9707 => "01110001",
 9708 => "10111101",
 9709 => "00000110",
 9710 => "11011110",
 9711 => "11101010",
 9712 => "10100100",
 9713 => "00100100",
 9714 => "00010011",
 9715 => "00100110",
 9716 => "11100010",
 9717 => "10100000",
 9718 => "00000001",
 9719 => "00010110",
 9720 => "10010111",
 9721 => "00110000",
 9722 => "01100000",
 9723 => "11110011",
 9724 => "01010110",
 9725 => "01100110",
 9726 => "01011100",
 9727 => "00010111",
 9728 => "10010111",
 9729 => "01100010",
 9730 => "10011011",
 9731 => "00000111",
 9732 => "00101010",
 9733 => "10010011",
 9734 => "01011111",
 9735 => "00101101",
 9736 => "10110000",
 9737 => "10110011",
 9738 => "01110111",
 9739 => "10001100",
 9740 => "11010001",
 9741 => "01001011",
 9742 => "00111000",
 9743 => "00010101",
 9744 => "11100110",
 9745 => "11100001",
 9746 => "11100010",
 9747 => "01000110",
 9748 => "10011000",
 9749 => "00101010",
 9750 => "10110101",
 9751 => "00110000",
 9752 => "00011110",
 9753 => "10011111",
 9754 => "11110001",
 9755 => "00000000",
 9756 => "01001111",
 9757 => "11000100",
 9758 => "00101101",
 9759 => "00110000",
 9760 => "11110000",
 9761 => "01010010",
 9762 => "01110011",
 9763 => "00100010",
 9764 => "01000011",
 9765 => "11101001",
 9766 => "11010010",
 9767 => "01001111",
 9768 => "11111011",
 9769 => "11000011",
 9770 => "00010011",
 9771 => "01100010",
 9772 => "11111011",
 9773 => "11110111",
 9774 => "10011011",
 9775 => "01011101",
 9776 => "00011111",
 9777 => "10101101",
 9778 => "10100010",
 9779 => "01001101",
 9780 => "00101110",
 9781 => "01111101",
 9782 => "01001101",
 9783 => "11101011",
 9784 => "00110011",
 9785 => "01001100",
 9786 => "11010110",
 9787 => "01100010",
 9788 => "01011100",
 9789 => "11111001",
 9790 => "00001000",
 9791 => "00101100",
 9792 => "01110010",
 9793 => "11001101",
 9794 => "10101110",
 9795 => "01010000",
 9796 => "10110100",
 9797 => "00110001",
 9798 => "00101010",
 9799 => "01111011",
 9800 => "11011011",
 9801 => "10001001",
 9802 => "00010001",
 9803 => "01101000",
 9804 => "01111100",
 9805 => "00001010",
 9806 => "00101011",
 9807 => "01111000",
 9808 => "00000010",
 9809 => "00010110",
 9810 => "10110011",
 9811 => "00011010",
 9812 => "11100010",
 9813 => "10010100",
 9814 => "11110111",
 9815 => "11111100",
 9816 => "10100100",
 9817 => "01101101",
 9818 => "10100000",
 9819 => "00000010",
 9820 => "10111110",
 9821 => "00110110",
 9822 => "01100001",
 9823 => "01110101",
 9824 => "00100010",
 9825 => "00100101",
 9826 => "11000100",
 9827 => "11010010",
 9828 => "10000110",
 9829 => "10101101",
 9830 => "01011100",
 9831 => "01001111",
 9832 => "00010000",
 9833 => "11110010",
 9834 => "11001101",
 9835 => "00011101",
 9836 => "01010000",
 9837 => "10101110",
 9838 => "10000101",
 9839 => "11000001",
 9840 => "11100100",
 9841 => "00100111",
 9842 => "10101100",
 9843 => "11001001",
 9844 => "01010110",
 9845 => "01111110",
 9846 => "01110011",
 9847 => "11000100",
 9848 => "11111100",
 9849 => "10111010",
 9850 => "11000000",
 9851 => "11111100",
 9852 => "11101100",
 9853 => "11110001",
 9854 => "11111110",
 9855 => "11100101",
 9856 => "00110110",
 9857 => "00110100",
 9858 => "10100110",
 9859 => "01111101",
 9860 => "11111011",
 9861 => "00011110",
 9862 => "01110100",
 9863 => "00100011",
 9864 => "00111011",
 9865 => "01101011",
 9866 => "01111100",
 9867 => "01010110",
 9868 => "11001011",
 9869 => "01001011",
 9870 => "00001010",
 9871 => "11100010",
 9872 => "10000011",
 9873 => "10010000",
 9874 => "11010010",
 9875 => "10111100",
 9876 => "01000000",
 9877 => "10001010",
 9878 => "00000110",
 9879 => "11011001",
 9880 => "00100010",
 9881 => "00110101",
 9882 => "01000100",
 9883 => "00110110",
 9884 => "10111111",
 9885 => "00011011",
 9886 => "00001110",
 9887 => "01101100",
 9888 => "01110001",
 9889 => "01000110",
 9890 => "10111100",
 9891 => "01100111",
 9892 => "01000000",
 9893 => "11001100",
 9894 => "11100110",
 9895 => "01100101",
 9896 => "01001101",
 9897 => "10101111",
 9898 => "01100011",
 9899 => "10011111",
 9900 => "01110101",
 9901 => "01000101",
 9902 => "10001001",
 9903 => "11101001",
 9904 => "01110101",
 9905 => "01101001",
 9906 => "00100000",
 9907 => "01010110",
 9908 => "01010101",
 9909 => "10100100",
 9910 => "01011010",
 9911 => "00110011",
 9912 => "01000101",
 9913 => "01011100",
 9914 => "11101110",
 9915 => "10111101",
 9916 => "01011111",
 9917 => "01000010",
 9918 => "01100101",
 9919 => "00101111",
 9920 => "11010100",
 9921 => "00000111",
 9922 => "00011011",
 9923 => "01010101",
 9924 => "11011001",
 9925 => "01001000",
 9926 => "00001010",
 9927 => "10000010",
 9928 => "01011001",
 9929 => "00000010",
 9930 => "00111001",
 9931 => "00110010",
 9932 => "11111010",
 9933 => "01000110",
 9934 => "00000000",
 9935 => "01001111",
 9936 => "10111010",
 9937 => "10111110",
 9938 => "10011010",
 9939 => "11010111",
 9940 => "00100011",
 9941 => "00101101",
 9942 => "00101100",
 9943 => "00101100",
 9944 => "00101011",
 9945 => "10001001",
 9946 => "11000000",
 9947 => "01001011",
 9948 => "01011011",
 9949 => "01111100",
 9950 => "01000011",
 9951 => "11100011",
 9952 => "11111001",
 9953 => "11001101",
 9954 => "11001100",
 9955 => "10000010",
 9956 => "11100100",
 9957 => "01010011",
 9958 => "10110001",
 9959 => "01001010",
 9960 => "01001101",
 9961 => "00011100",
 9962 => "10011000",
 9963 => "11001011",
 9964 => "00100000",
 9965 => "11110100",
 9966 => "01110000",
 9967 => "00100101",
 9968 => "11110011",
 9969 => "00101010",
 9970 => "10100000",
 9971 => "10100111",
 9972 => "00110001",
 9973 => "11000001",
 9974 => "11110010",
 9975 => "10010001",
 9976 => "01000011",
 9977 => "10101001",
 9978 => "10001000",
 9979 => "10111110",
 9980 => "00100101",
 9981 => "01111000",
 9982 => "00000000",
 9983 => "00101010",
 9984 => "00100110",
 9985 => "10100101",
 9986 => "10001000",
 9987 => "10010000",
 9988 => "10000101",
 9989 => "00110001",
 9990 => "01001101",
 9991 => "10000001",
 9992 => "01011110",
 9993 => "00010000",
 9994 => "10011001",
 9995 => "11011001",
 9996 => "00011011",
 9997 => "10010101",
 9998 => "01110100",
 9999 => "11010101",
 10000 => "11100101",
 10001 => "10000111",
 10002 => "00010000",
 10003 => "00101001",
 10004 => "10011011",
 10005 => "01110011",
 10006 => "01101100",
 10007 => "10100111",
 10008 => "11011000",
 10009 => "10001110",
 10010 => "01110111",
 10011 => "10010001",
 10012 => "10001110",
 10013 => "10101001",
 10014 => "00010101",
 10015 => "11011010",
 10016 => "11010010",
 10017 => "00111000",
 10018 => "10101100",
 10019 => "00010001",
 10020 => "11111101",
 10021 => "01100010",
 10022 => "11011101",
 10023 => "10001010",
 10024 => "00000110",
 10025 => "01111110",
 10026 => "11001011",
 10027 => "01111111",
 10028 => "01101110",
 10029 => "01100101",
 10030 => "11011100",
 10031 => "11101101",
 10032 => "00111000",
 10033 => "11000011",
 10034 => "01011001",
 10035 => "10100011",
 10036 => "00011111",
 10037 => "10111111",
 10038 => "11110010",
 10039 => "11001100",
 10040 => "10111011",
 10041 => "00010011",
 10042 => "01001101",
 10043 => "10000001",
 10044 => "11101011",
 10045 => "00111000",
 10046 => "10100110",
 10047 => "00111011",
 10048 => "10011010",
 10049 => "01001111",
 10050 => "10100101",
 10051 => "00101111",
 10052 => "00010011",
 10053 => "00010010",
 10054 => "00101010",
 10055 => "10010101",
 10056 => "10111010",
 10057 => "01011111",
 10058 => "01000010",
 10059 => "10111011",
 10060 => "00000111",
 10061 => "00010111",
 10062 => "10011000",
 10063 => "00000011",
 10064 => "10110011",
 10065 => "00000011",
 10066 => "01100111",
 10067 => "11101001",
 10068 => "10010110",
 10069 => "11100111",
 10070 => "11101111",
 10071 => "11000100",
 10072 => "01111101",
 10073 => "11000100",
 10074 => "00000011",
 10075 => "01010000",
 10076 => "11010111",
 10077 => "11000111",
 10078 => "00010100",
 10079 => "01011111",
 10080 => "01010001",
 10081 => "11111001",
 10082 => "00100011",
 10083 => "10010111",
 10084 => "11010111",
 10085 => "01010111",
 10086 => "11011010",
 10087 => "11101110",
 10088 => "00100101",
 10089 => "00001100",
 10090 => "11110001",
 10091 => "00001100",
 10092 => "11001111",
 10093 => "01000001",
 10094 => "11010000",
 10095 => "11000100",
 10096 => "10011010",
 10097 => "11010010",
 10098 => "01001110",
 10099 => "10100001",
 10100 => "11001110",
 10101 => "00011000",
 10102 => "11111000",
 10103 => "00110111",
 10104 => "10010000",
 10105 => "00010010",
 10106 => "11101001",
 10107 => "00011100",
 10108 => "00110011",
 10109 => "00101011",
 10110 => "01000111",
 10111 => "01100110",
 10112 => "11100010",
 10113 => "01100010",
 10114 => "11101100",
 10115 => "00011011",
 10116 => "00101111",
 10117 => "10011011",
 10118 => "00101000",
 10119 => "10111110",
 10120 => "10011010",
 10121 => "01110110",
 10122 => "00010111",
 10123 => "00010110",
 10124 => "10101011",
 10125 => "01110010",
 10126 => "10111110",
 10127 => "00000000",
 10128 => "00101110",
 10129 => "00001110",
 10130 => "10100011",
 10131 => "11010010",
 10132 => "10111110",
 10133 => "01000110",
 10134 => "11011101",
 10135 => "01100001",
 10136 => "10110100",
 10137 => "00111100",
 10138 => "10011010",
 10139 => "00011000",
 10140 => "01010100",
 10141 => "01000111",
 10142 => "00000011",
 10143 => "01000101",
 10144 => "10101110",
 10145 => "01111100",
 10146 => "01101010",
 10147 => "01011000",
 10148 => "01100110",
 10149 => "11011010",
 10150 => "11011001",
 10151 => "01101001",
 10152 => "11000011",
 10153 => "11111100",
 10154 => "10001111",
 10155 => "11000010",
 10156 => "00110111",
 10157 => "01111000",
 10158 => "10110000",
 10159 => "10110100",
 10160 => "00101110",
 10161 => "00000100",
 10162 => "10111101",
 10163 => "01101010",
 10164 => "01101000",
 10165 => "01000111",
 10166 => "10111100",
 10167 => "10010101",
 10168 => "10001001",
 10169 => "00010110",
 10170 => "01101010",
 10171 => "01101110",
 10172 => "10000101",
 10173 => "11100101",
 10174 => "00100110",
 10175 => "10011101",
 10176 => "11000111",
 10177 => "10111001",
 10178 => "01001011",
 10179 => "01110100",
 10180 => "00110011",
 10181 => "00010111",
 10182 => "01100011",
 10183 => "01101110",
 10184 => "00111101",
 10185 => "00010101",
 10186 => "01011011",
 10187 => "10001111",
 10188 => "11110010",
 10189 => "00000110",
 10190 => "11000111",
 10191 => "01111111",
 10192 => "01111011",
 10193 => "11010000",
 10194 => "11101001",
 10195 => "10010001",
 10196 => "10111001",
 10197 => "01011110",
 10198 => "01010000",
 10199 => "01010010",
 10200 => "00110000",
 10201 => "11111101",
 10202 => "10011101",
 10203 => "01000111",
 10204 => "00010101",
 10205 => "00011011",
 10206 => "00011001",
 10207 => "10011111",
 10208 => "01101010",
 10209 => "00101011",
 10210 => "01101101",
 10211 => "10111111",
 10212 => "11011000",
 10213 => "10110101",
 10214 => "11111001",
 10215 => "10111001",
 10216 => "01001011",
 10217 => "00100010",
 10218 => "11001001",
 10219 => "10000011",
 10220 => "11100001",
 10221 => "00111010",
 10222 => "10011100",
 10223 => "00011110",
 10224 => "11101010",
 10225 => "10011100",
 10226 => "01010100",
 10227 => "01000110",
 10228 => "11101111",
 10229 => "11001101",
 10230 => "00110001",
 10231 => "10001110",
 10232 => "11100100",
 10233 => "00000011",
 10234 => "10101011",
 10235 => "00010111",
 10236 => "00011000",
 10237 => "11111001",
 10238 => "10010111",
 10239 => "01111110",
 10240 => "10011011",
 10241 => "01100000",
 10242 => "10110110",
 10243 => "10101010",
 10244 => "00001001",
 10245 => "01111100",
 10246 => "11111010",
 10247 => "00001111",
 10248 => "10000001",
 10249 => "10001100",
 10250 => "00011110",
 10251 => "11001010",
 10252 => "10001000",
 10253 => "01111101",
 10254 => "00001000",
 10255 => "01100011",
 10256 => "11111001",
 10257 => "01100101",
 10258 => "00011110",
 10259 => "01111110",
 10260 => "01101001",
 10261 => "01110011",
 10262 => "10000110",
 10263 => "00111000",
 10264 => "10011000",
 10265 => "01101000",
 10266 => "11001110",
 10267 => "10100100",
 10268 => "10100101",
 10269 => "10001111",
 10270 => "11100101",
 10271 => "00110011",
 10272 => "11011100",
 10273 => "11011000",
 10274 => "00101011",
 10275 => "01001100",
 10276 => "10011101",
 10277 => "01101000",
 10278 => "01111100",
 10279 => "00101100",
 10280 => "10001111",
 10281 => "11011011",
 10282 => "11011111",
 10283 => "10000111",
 10284 => "10111100",
 10285 => "10110111",
 10286 => "11100010",
 10287 => "10101100",
 10288 => "00011100",
 10289 => "11011101",
 10290 => "11011000",
 10291 => "00000000",
 10292 => "01100010",
 10293 => "00110100",
 10294 => "11111100",
 10295 => "00010000",
 10296 => "11001011",
 10297 => "01000000",
 10298 => "10011100",
 10299 => "11100001",
 10300 => "10110101",
 10301 => "01110100",
 10302 => "11111101",
 10303 => "11001010",
 10304 => "10010101",
 10305 => "11111101",
 10306 => "10111001",
 10307 => "01010001",
 10308 => "11101010",
 10309 => "10100101",
 10310 => "00110011",
 10311 => "11011101",
 10312 => "10111001",
 10313 => "01101010",
 10314 => "00000100",
 10315 => "00110110",
 10316 => "10100010",
 10317 => "01100111",
 10318 => "01110101",
 10319 => "00101011",
 10320 => "01111111",
 10321 => "00111100",
 10322 => "11001001",
 10323 => "10000001",
 10324 => "00100001",
 10325 => "11110000",
 10326 => "11110101",
 10327 => "01110010",
 10328 => "01111100",
 10329 => "10000101",
 10330 => "11110110",
 10331 => "10000011",
 10332 => "11100111",
 10333 => "00001110",
 10334 => "01010001",
 10335 => "01000110",
 10336 => "01111111",
 10337 => "00100010",
 10338 => "01100011",
 10339 => "01111010",
 10340 => "10100100",
 10341 => "11000100",
 10342 => "01111110",
 10343 => "11100011",
 10344 => "11001000",
 10345 => "01011110",
 10346 => "10110000",
 10347 => "10100000",
 10348 => "00000011",
 10349 => "01000111",
 10350 => "10001011",
 10351 => "10100001",
 10352 => "11100110",
 10353 => "11001011",
 10354 => "01101100",
 10355 => "00100111",
 10356 => "10000100",
 10357 => "10100011",
 10358 => "11000011",
 10359 => "11100011",
 10360 => "00110000",
 10361 => "00110001",
 10362 => "10100110",
 10363 => "00011011",
 10364 => "01111001",
 10365 => "00100011",
 10366 => "11100111",
 10367 => "10101101",
 10368 => "11100100",
 10369 => "11010010",
 10370 => "11111000",
 10371 => "11010101",
 10372 => "11011001",
 10373 => "00011010",
 10374 => "01101001",
 10375 => "01000011",
 10376 => "11101000",
 10377 => "11011001",
 10378 => "10111110",
 10379 => "01000001",
 10380 => "10000001",
 10381 => "00111101",
 10382 => "01111001",
 10383 => "01101100",
 10384 => "01111100",
 10385 => "00111111",
 10386 => "10100111",
 10387 => "10110000",
 10388 => "00000111",
 10389 => "01111100",
 10390 => "00111111",
 10391 => "00101101",
 10392 => "10010001",
 10393 => "11100000",
 10394 => "01001000",
 10395 => "11000000",
 10396 => "00011100",
 10397 => "11010100",
 10398 => "10100010",
 10399 => "00001000",
 10400 => "01000011",
 10401 => "11010110",
 10402 => "01011100",
 10403 => "10010111",
 10404 => "00001111",
 10405 => "10000010",
 10406 => "11100101",
 10407 => "00111111",
 10408 => "00001010",
 10409 => "11000001",
 10410 => "11111010",
 10411 => "11101011",
 10412 => "11101000",
 10413 => "10000111",
 10414 => "11100100",
 10415 => "01011001",
 10416 => "11011110",
 10417 => "01000101",
 10418 => "11100110",
 10419 => "11101001",
 10420 => "00101001",
 10421 => "01001011",
 10422 => "10010010",
 10423 => "00100100",
 10424 => "00011101",
 10425 => "00011000",
 10426 => "10001000",
 10427 => "00011101",
 10428 => "10110011",
 10429 => "00010010",
 10430 => "01000011",
 10431 => "11011000",
 10432 => "11110011",
 10433 => "11001011",
 10434 => "00111011",
 10435 => "11001001",
 10436 => "01101100",
 10437 => "10101000",
 10438 => "01101011",
 10439 => "01110010",
 10440 => "10111010",
 10441 => "01100000",
 10442 => "00000001",
 10443 => "10010110",
 10444 => "11001111",
 10445 => "10001000",
 10446 => "01100111",
 10447 => "01111001",
 10448 => "01111101",
 10449 => "00101000",
 10450 => "11111010",
 10451 => "01110000",
 10452 => "01010111",
 10453 => "11101011",
 10454 => "10110000",
 10455 => "11101011",
 10456 => "10110011",
 10457 => "00000001",
 10458 => "00110011",
 10459 => "11101000",
 10460 => "11110000",
 10461 => "11000011",
 10462 => "10110001",
 10463 => "10111110",
 10464 => "10111110",
 10465 => "10011000",
 10466 => "00000000",
 10467 => "11100001",
 10468 => "00101001",
 10469 => "10101011",
 10470 => "00111101",
 10471 => "00011001",
 10472 => "00010000",
 10473 => "11101000",
 10474 => "10111110",
 10475 => "10001010",
 10476 => "01010111",
 10477 => "00001001",
 10478 => "11111011",
 10479 => "00001100",
 10480 => "01101101",
 10481 => "00000010",
 10482 => "01101011",
 10483 => "10011100",
 10484 => "11010011",
 10485 => "11011001",
 10486 => "00100110",
 10487 => "11101100",
 10488 => "10111111",
 10489 => "10110100",
 10490 => "11000001",
 10491 => "10011000",
 10492 => "11100110",
 10493 => "00110111",
 10494 => "01101000",
 10495 => "10100101",
 10496 => "10000100",
 10497 => "11010000",
 10498 => "00101011",
 10499 => "11101101",
 10500 => "00110101",
 10501 => "11001000",
 10502 => "10101100",
 10503 => "10111001",
 10504 => "10011000",
 10505 => "00100001",
 10506 => "10001111",
 10507 => "10011111",
 10508 => "10100100",
 10509 => "01101111",
 10510 => "01001100",
 10511 => "11100000",
 10512 => "11110100",
 10513 => "01001111",
 10514 => "10000011",
 10515 => "00010011",
 10516 => "00010011",
 10517 => "10110001",
 10518 => "01101001",
 10519 => "01100110",
 10520 => "01010111",
 10521 => "01110000",
 10522 => "00100001",
 10523 => "10111011",
 10524 => "10010100",
 10525 => "11011011",
 10526 => "00010011",
 10527 => "10010110",
 10528 => "10011010",
 10529 => "00010111",
 10530 => "00101111",
 10531 => "01111001",
 10532 => "01000011",
 10533 => "10100111",
 10534 => "01100000",
 10535 => "11111010",
 10536 => "11001010",
 10537 => "01010100",
 10538 => "10111111",
 10539 => "01001011",
 10540 => "11111001",
 10541 => "11001000",
 10542 => "10110010",
 10543 => "11000101",
 10544 => "10011011",
 10545 => "00010011",
 10546 => "11000010",
 10547 => "00011101",
 10548 => "11011011",
 10549 => "10101010",
 10550 => "00110001",
 10551 => "10011001",
 10552 => "01111000",
 10553 => "00101001",
 10554 => "01001010",
 10555 => "01110001",
 10556 => "11011110",
 10557 => "01011010",
 10558 => "01100101",
 10559 => "10011101",
 10560 => "11111110",
 10561 => "10110001",
 10562 => "10010011",
 10563 => "00100001",
 10564 => "00101111",
 10565 => "01011010",
 10566 => "10001111",
 10567 => "11001000",
 10568 => "11000101",
 10569 => "00001101",
 10570 => "01100110",
 10571 => "01101101",
 10572 => "10100011",
 10573 => "10010111",
 10574 => "01100011",
 10575 => "10100101",
 10576 => "11010001",
 10577 => "01011111",
 10578 => "01011110",
 10579 => "11001001",
 10580 => "11110010",
 10581 => "00111001",
 10582 => "10011100",
 10583 => "01111011",
 10584 => "01110011",
 10585 => "00010110",
 10586 => "11001001",
 10587 => "10101100",
 10588 => "00010011",
 10589 => "01101000",
 10590 => "10000110",
 10591 => "00101101",
 10592 => "01011100",
 10593 => "00000000",
 10594 => "00010010",
 10595 => "10011001",
 10596 => "00000000",
 10597 => "00010011",
 10598 => "00100000",
 10599 => "10010010",
 10600 => "11100110",
 10601 => "01001011",
 10602 => "01100110",
 10603 => "11010001",
 10604 => "10100011",
 10605 => "11000001",
 10606 => "00100011",
 10607 => "01100101",
 10608 => "10011110",
 10609 => "11000001",
 10610 => "00010101",
 10611 => "00111010",
 10612 => "01110100",
 10613 => "00111111",
 10614 => "11111100",
 10615 => "10101010",
 10616 => "01100000",
 10617 => "10000010",
 10618 => "01100011",
 10619 => "00110101",
 10620 => "01101111",
 10621 => "01111001",
 10622 => "11011111",
 10623 => "10000100",
 10624 => "10111100",
 10625 => "10111000",
 10626 => "11011111",
 10627 => "11101110",
 10628 => "01010000",
 10629 => "11111111",
 10630 => "00001101",
 10631 => "10011000",
 10632 => "00111011",
 10633 => "01101111",
 10634 => "11100100",
 10635 => "11000101",
 10636 => "11110110",
 10637 => "10101000",
 10638 => "10100111",
 10639 => "10110110",
 10640 => "01100011",
 10641 => "01100010",
 10642 => "10001101",
 10643 => "10011001",
 10644 => "10011111",
 10645 => "00111001",
 10646 => "10011011",
 10647 => "01001000",
 10648 => "10110010",
 10649 => "01111101",
 10650 => "00000011",
 10651 => "01000010",
 10652 => "01001001",
 10653 => "10100100",
 10654 => "10110010",
 10655 => "00000111",
 10656 => "01110001",
 10657 => "01010000",
 10658 => "11000110",
 10659 => "01011101",
 10660 => "01110010",
 10661 => "00100000",
 10662 => "11110000",
 10663 => "00111111",
 10664 => "11001101",
 10665 => "00011100",
 10666 => "01110101",
 10667 => "01011000",
 10668 => "00011111",
 10669 => "00100000",
 10670 => "10100110",
 10671 => "11100101",
 10672 => "10010100",
 10673 => "01111010",
 10674 => "11100001",
 10675 => "10101010",
 10676 => "00001001",
 10677 => "11010000",
 10678 => "00011101",
 10679 => "11000100",
 10680 => "01011110",
 10681 => "11110100",
 10682 => "01101110",
 10683 => "11111111",
 10684 => "00100111",
 10685 => "10001000",
 10686 => "11010110",
 10687 => "11011110",
 10688 => "10000110",
 10689 => "11101110",
 10690 => "01101100",
 10691 => "11001111",
 10692 => "11101111",
 10693 => "10000110",
 10694 => "10010100",
 10695 => "00011110",
 10696 => "00000000",
 10697 => "01110011",
 10698 => "01101001",
 10699 => "01111101",
 10700 => "00010111",
 10701 => "10101001",
 10702 => "00111010",
 10703 => "10010100",
 10704 => "11000100",
 10705 => "10110011",
 10706 => "01110011",
 10707 => "10000111",
 10708 => "01000101",
 10709 => "10110000",
 10710 => "00111111",
 10711 => "11111110",
 10712 => "01100100",
 10713 => "00100100",
 10714 => "10111010",
 10715 => "10110010",
 10716 => "00010111",
 10717 => "01011100",
 10718 => "00111101",
 10719 => "00010110",
 10720 => "00100010",
 10721 => "11011101",
 10722 => "11110010",
 10723 => "00100011",
 10724 => "11100101",
 10725 => "10111001",
 10726 => "00111000",
 10727 => "11010100",
 10728 => "00010101",
 10729 => "01001000",
 10730 => "11000001",
 10731 => "11110111",
 10732 => "00111100",
 10733 => "11100011",
 10734 => "01111110",
 10735 => "10111100",
 10736 => "11011001",
 10737 => "01011010",
 10738 => "10100110",
 10739 => "00110011",
 10740 => "01001011",
 10741 => "11100101",
 10742 => "01100010",
 10743 => "01010000",
 10744 => "01001000",
 10745 => "01001001",
 10746 => "10000110",
 10747 => "10011000",
 10748 => "11011011",
 10749 => "00010001",
 10750 => "11011011",
 10751 => "11101010",
 10752 => "10011001",
 10753 => "10010000",
 10754 => "10101110",
 10755 => "00000100",
 10756 => "01111000",
 10757 => "10000010",
 10758 => "01010111",
 10759 => "10001001",
 10760 => "10100001",
 10761 => "00000101",
 10762 => "00101101",
 10763 => "10110001",
 10764 => "11011011",
 10765 => "01010000",
 10766 => "11011111",
 10767 => "10100000",
 10768 => "11000000",
 10769 => "01010111",
 10770 => "10000010",
 10771 => "01000101",
 10772 => "10011000",
 10773 => "10001101",
 10774 => "01110010",
 10775 => "11011101",
 10776 => "01110110",
 10777 => "01010000",
 10778 => "01111001",
 10779 => "01100000",
 10780 => "00101011",
 10781 => "10010010",
 10782 => "10000100",
 10783 => "01011000",
 10784 => "01111010",
 10785 => "00100111",
 10786 => "10101100",
 10787 => "00111010",
 10788 => "10101011",
 10789 => "00001001",
 10790 => "00010100",
 10791 => "10110111",
 10792 => "01001101",
 10793 => "00000001",
 10794 => "01001000",
 10795 => "01110101",
 10796 => "01000011",
 10797 => "00000101",
 10798 => "11001011",
 10799 => "11111011",
 10800 => "01010001",
 10801 => "00101110",
 10802 => "01101111",
 10803 => "10000010",
 10804 => "00000001",
 10805 => "01100001",
 10806 => "01100011",
 10807 => "01000101",
 10808 => "11110111",
 10809 => "11001001",
 10810 => "10000010",
 10811 => "01000011",
 10812 => "00010000",
 10813 => "11111000",
 10814 => "11110001",
 10815 => "11100100",
 10816 => "00001000",
 10817 => "10100001",
 10818 => "11110010",
 10819 => "10111101",
 10820 => "01111000",
 10821 => "11110101",
 10822 => "10100011",
 10823 => "11011111",
 10824 => "00111111",
 10825 => "01001000",
 10826 => "01111111",
 10827 => "01110001",
 10828 => "10111000",
 10829 => "00001101",
 10830 => "01110010",
 10831 => "01001110",
 10832 => "00101011",
 10833 => "11001110",
 10834 => "10010010",
 10835 => "00010100",
 10836 => "11001111",
 10837 => "01110011",
 10838 => "11001101",
 10839 => "00001100",
 10840 => "11111100",
 10841 => "11100101",
 10842 => "00110111",
 10843 => "01011010",
 10844 => "01100000",
 10845 => "00010000",
 10846 => "10111110",
 10847 => "11000110",
 10848 => "01001011",
 10849 => "00110001",
 10850 => "11111011",
 10851 => "01000100",
 10852 => "00101001",
 10853 => "10010001",
 10854 => "00000011",
 10855 => "01100111",
 10856 => "00101111",
 10857 => "01101000",
 10858 => "11101000",
 10859 => "11100010",
 10860 => "10010011",
 10861 => "00000111",
 10862 => "00110000",
 10863 => "00010011",
 10864 => "11010011",
 10865 => "10001001",
 10866 => "00100010",
 10867 => "01001001",
 10868 => "10101010",
 10869 => "11100101",
 10870 => "10101001",
 10871 => "01111110",
 10872 => "10110110",
 10873 => "01110011",
 10874 => "01000001",
 10875 => "10011000",
 10876 => "10110011",
 10877 => "00111100",
 10878 => "01010100",
 10879 => "00100011",
 10880 => "11110101",
 10881 => "01101101",
 10882 => "11001110",
 10883 => "10111001",
 10884 => "11111110",
 10885 => "01011111",
 10886 => "10000001",
 10887 => "00011001",
 10888 => "01011110",
 10889 => "01111000",
 10890 => "00000001",
 10891 => "11001001",
 10892 => "01101110",
 10893 => "10010111",
 10894 => "11101101",
 10895 => "00011111",
 10896 => "01110111",
 10897 => "10101111",
 10898 => "10001101",
 10899 => "01001110",
 10900 => "10010001",
 10901 => "10111001",
 10902 => "00010101",
 10903 => "01001110",
 10904 => "11000001",
 10905 => "10011010",
 10906 => "00010010", others => (others =>'0'));
component project_reti_logiche is 
    port (
            i_clk         : in  std_logic;
            i_start       : in  std_logic;
            i_rst         : in  std_logic;
            i_data       : in  std_logic_vector(7 downto 0); --1 byte
            o_address     : out std_logic_vector(15 downto 0); --16 bit addr: max size is 255*255 + 3 more for max x and y and thresh.
            o_done            : out std_logic;
            o_en         : out std_logic;
            o_we       : out std_logic;
            o_data            : out std_logic_vector (7 downto 0)
          );
end component project_reti_logiche;
begin 
	UUT: project_reti_logiche
	port map (
		  i_clk      	=> tb_clk,	
          i_start       => tb_start,
          i_rst      	=> tb_rst,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address, 
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
		  o_we 	=> mem_we,
          o_data    => mem_i_data
);p_CLK_GEN : process is
  begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
  end process p_CLK_GEN; 
 MEM : process(tb_clk)
   begin
    if tb_clk'event and tb_clk = '1' then
     if enable_wire = '1' then
      if mem_we = '1' then
       RAM(conv_integer(mem_address))              <= mem_i_data;
       mem_o_data                      <= mem_i_data;
      else
       mem_o_data <= RAM(conv_integer(mem_address));
      end if;
     end if;
    end if;
   end process;
test : process is
begin 
wait for 100 ns;
wait for c_CLOCK_PERIOD;
tb_rst <= '1';
wait for c_CLOCK_PERIOD;
tb_rst <= '0';
wait for c_CLOCK_PERIOD;
tb_start <= '1';
wait for c_CLOCK_PERIOD; 
tb_start <= '0';
wait until tb_done = '1';
wait until tb_done = '0';
wait until rising_edge(tb_clk);

 
assert RAM(1) = "00101010" report "FAIL high bits" severity failure;
assert RAM(0) = "10010110" report "FAIL low bits" severity failure;
assert false report "Simulation Ended!, test passed" severity failure;
end process test;
 end projecttb;